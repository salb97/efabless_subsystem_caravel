VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbytes_1rw1r_200x48_8
   CLASS BLOCK ;
   SIZE 1532.42 BY 349.9 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  352.92 0.0 353.3 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  358.36 0.0 358.74 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  364.48 0.0 364.86 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  370.6 0.0 370.98 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  376.04 0.0 376.42 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  382.16 0.0 382.54 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  386.92 0.0 387.3 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  393.72 0.0 394.1 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  399.16 0.0 399.54 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 404.98 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  411.4 0.0 411.78 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  416.16 0.0 416.54 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  422.96 0.0 423.34 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  429.08 0.0 429.46 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  434.52 0.0 434.9 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  439.96 0.0 440.34 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  445.4 0.0 445.78 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  452.2 0.0 452.58 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  457.64 0.0 458.02 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  463.76 0.0 464.14 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  468.52 0.0 468.9 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  475.32 0.0 475.7 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  480.76 0.0 481.14 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  486.88 0.0 487.26 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 0.0 492.7 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  497.76 0.0 498.14 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  503.88 0.0 504.26 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  510.68 0.0 511.06 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  515.44 0.0 515.82 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  521.56 0.0 521.94 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  527.68 0.0 528.06 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  533.12 0.0 533.5 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  539.24 0.0 539.62 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  544.68 0.0 545.06 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  550.8 0.0 551.18 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  556.24 0.0 556.62 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  562.36 0.0 562.74 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  569.16 0.0 569.54 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  573.92 0.0 574.3 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  580.72 0.0 581.1 1.06 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  585.48 0.0 585.86 1.06 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  592.28 0.0 592.66 1.06 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  597.72 0.0 598.1 1.06 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  603.84 0.0 604.22 1.06 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  609.28 0.0 609.66 1.06 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  615.4 0.0 615.78 1.06 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  620.84 0.0 621.22 1.06 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  626.96 0.0 627.34 1.06 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  632.4 0.0 632.78 1.06 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  639.2 0.0 639.58 1.06 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  643.96 0.0 644.34 1.06 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  650.76 0.0 651.14 1.06 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  656.2 0.0 656.58 1.06 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  662.32 0.0 662.7 1.06 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  668.44 0.0 668.82 1.06 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  673.88 0.0 674.26 1.06 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  680.0 0.0 680.38 1.06 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  684.76 0.0 685.14 1.06 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  691.56 0.0 691.94 1.06 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  696.32 0.0 696.7 1.06 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  702.44 0.0 702.82 1.06 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  709.24 0.0 709.62 1.06 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  714.0 0.0 714.38 1.06 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  720.8 0.0 721.18 1.06 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  726.92 0.0 727.3 1.06 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  732.36 0.0 732.74 1.06 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  738.48 0.0 738.86 1.06 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  743.24 0.0 743.62 1.06 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  749.36 0.0 749.74 1.06 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  754.8 0.0 755.18 1.06 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  760.92 0.0 761.3 1.06 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  766.36 0.0 766.74 1.06 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  772.48 0.0 772.86 1.06 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  778.6 0.0 778.98 1.06 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  784.04 0.0 784.42 1.06 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  790.16 0.0 790.54 1.06 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  796.28 0.0 796.66 1.06 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  802.4 0.0 802.78 1.06 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  808.52 0.0 808.9 1.06 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  813.96 0.0 814.34 1.06 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  820.08 0.0 820.46 1.06 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  825.52 0.0 825.9 1.06 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  831.64 0.0 832.02 1.06 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  837.08 0.0 837.46 1.06 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  842.52 0.0 842.9 1.06 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  849.32 0.0 849.7 1.06 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  854.08 0.0 854.46 1.06 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  860.88 0.0 861.26 1.06 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  865.64 0.0 866.02 1.06 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  872.44 0.0 872.82 1.06 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  878.56 0.0 878.94 1.06 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  884.0 0.0 884.38 1.06 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  889.44 0.0 889.82 1.06 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  894.88 0.0 895.26 1.06 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  901.0 0.0 901.38 1.06 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  907.12 0.0 907.5 1.06 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  912.56 0.0 912.94 1.06 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  918.68 0.0 919.06 1.06 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  924.12 0.0 924.5 1.06 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  930.92 0.0 931.3 1.06 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  937.04 0.0 937.42 1.06 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  941.8 0.0 942.18 1.06 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  947.92 0.0 948.3 1.06 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  953.36 0.0 953.74 1.06 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  959.48 0.0 959.86 1.06 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  965.6 0.0 965.98 1.06 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  971.04 0.0 971.42 1.06 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  977.84 0.0 978.22 1.06 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  982.6 0.0 982.98 1.06 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  989.4 0.0 989.78 1.06 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  994.84 0.0 995.22 1.06 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1000.96 0.0 1001.34 1.06 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1007.08 0.0 1007.46 1.06 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1011.84 0.0 1012.22 1.06 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1018.64 0.0 1019.02 1.06 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1023.4 0.0 1023.78 1.06 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1029.52 0.0 1029.9 1.06 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1036.32 0.0 1036.7 1.06 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1041.08 0.0 1041.46 1.06 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1047.88 0.0 1048.26 1.06 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1053.32 0.0 1053.7 1.06 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1059.44 0.0 1059.82 1.06 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1065.56 0.0 1065.94 1.06 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1070.32 0.0 1070.7 1.06 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1077.12 0.0 1077.5 1.06 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1082.56 0.0 1082.94 1.06 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1088.68 0.0 1089.06 1.06 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1094.12 0.0 1094.5 1.06 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1100.24 0.0 1100.62 1.06 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1105.68 0.0 1106.06 1.06 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1111.8 0.0 1112.18 1.06 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1117.24 0.0 1117.62 1.06 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1122.68 0.0 1123.06 1.06 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1128.8 0.0 1129.18 1.06 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1135.6 0.0 1135.98 1.06 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1140.36 0.0 1140.74 1.06 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1146.48 0.0 1146.86 1.06 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1152.6 0.0 1152.98 1.06 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1158.72 0.0 1159.1 1.06 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1163.48 0.0 1163.86 1.06 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1169.6 0.0 1169.98 1.06 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1175.72 0.0 1176.1 1.06 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1181.16 0.0 1181.54 1.06 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1187.28 0.0 1187.66 1.06 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1194.08 0.0 1194.46 1.06 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1198.84 0.0 1199.22 1.06 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1205.64 0.0 1206.02 1.06 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1210.4 0.0 1210.78 1.06 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1217.2 0.0 1217.58 1.06 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1223.32 0.0 1223.7 1.06 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1228.76 0.0 1229.14 1.06 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1234.2 0.0 1234.58 1.06 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1240.32 0.0 1240.7 1.06 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1245.76 0.0 1246.14 1.06 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1251.2 0.0 1251.58 1.06 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1257.32 0.0 1257.7 1.06 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1264.12 0.0 1264.5 1.06 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1269.56 0.0 1269.94 1.06 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1275.0 0.0 1275.38 1.06 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1281.12 0.0 1281.5 1.06 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1287.24 0.0 1287.62 1.06 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1292.0 0.0 1292.38 1.06 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1298.8 0.0 1299.18 1.06 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1304.24 0.0 1304.62 1.06 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1309.68 0.0 1310.06 1.06 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1315.8 0.0 1316.18 1.06 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1322.6 0.0 1322.98 1.06 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1327.36 0.0 1327.74 1.06 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1333.48 0.0 1333.86 1.06 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1338.92 0.0 1339.3 1.06 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1345.72 0.0 1346.1 1.06 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1350.48 0.0 1350.86 1.06 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1357.28 0.0 1357.66 1.06 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1362.04 0.0 1362.42 1.06 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1368.84 0.0 1369.22 1.06 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1374.28 0.0 1374.66 1.06 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1379.72 0.0 1380.1 1.06 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1385.84 0.0 1386.22 1.06 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1391.96 0.0 1392.34 1.06 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1397.4 0.0 1397.78 1.06 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1403.52 0.0 1403.9 1.06 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1408.96 0.0 1409.34 1.06 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1415.08 0.0 1415.46 1.06 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1421.88 0.0 1422.26 1.06 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1427.32 0.0 1427.7 1.06 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1433.44 0.0 1433.82 1.06 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1438.88 0.0 1439.26 1.06 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1445.0 0.0 1445.38 1.06 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1450.44 0.0 1450.82 1.06 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1456.56 0.0 1456.94 1.06 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1462.68 0.0 1463.06 1.06 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1467.44 0.0 1467.82 1.06 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1474.24 0.0 1474.62 1.06 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1479.0 0.0 1479.38 1.06 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1485.8 0.0 1486.18 1.06 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1490.56 0.0 1490.94 1.06 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1497.36 0.0 1497.74 1.06 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1503.48 0.0 1503.86 1.06 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1508.92 0.0 1509.3 1.06 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1514.36 0.0 1514.74 1.06 ;
      END
   END din0[199]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 348.84 197.58 349.9 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 348.84 192.82 349.9 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.52 348.84 196.9 349.9 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 348.84 193.5 349.9 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.84 348.84 196.22 349.9 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.16 348.84 195.54 349.9 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  966.96 348.84 967.34 349.9 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  967.64 348.84 968.02 349.9 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  966.28 348.84 966.66 349.9 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  966.28 0.0 966.66 1.06 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  967.64 0.0 968.02 1.06 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  966.96 0.0 967.34 1.06 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.68 1.06 137.06 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1147.84 348.84 1148.22 349.9 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 145.52 1.06 145.9 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 138.04 1.06 138.42 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1130.16 348.84 1130.54 349.9 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.72 0.0 207.1 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.16 0.0 212.54 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.72 0.0 224.1 1.06 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 0.0 230.9 1.06 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 1.06 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 1.06 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 0.0 247.9 1.06 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 0.0 254.02 1.06 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.08 0.0 259.46 1.06 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.52 0.0 264.9 1.06 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  271.32 0.0 271.7 1.06 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 1.06 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.2 0.0 282.58 1.06 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  287.64 0.0 288.02 1.06 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.76 0.0 294.14 1.06 ;
      END
   END wmask0[15]
   PIN wmask0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  299.2 0.0 299.58 1.06 ;
      END
   END wmask0[16]
   PIN wmask0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  305.32 0.0 305.7 1.06 ;
      END
   END wmask0[17]
   PIN wmask0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  312.12 0.0 312.5 1.06 ;
      END
   END wmask0[18]
   PIN wmask0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  316.88 0.0 317.26 1.06 ;
      END
   END wmask0[19]
   PIN wmask0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  323.68 0.0 324.06 1.06 ;
      END
   END wmask0[20]
   PIN wmask0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  329.12 0.0 329.5 1.06 ;
      END
   END wmask0[21]
   PIN wmask0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  334.56 0.0 334.94 1.06 ;
      END
   END wmask0[22]
   PIN wmask0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  340.68 0.0 341.06 1.06 ;
      END
   END wmask0[23]
   PIN wmask0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  346.12 0.0 346.5 1.06 ;
      END
   END wmask0[24]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 0.0 268.3 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  277.44 0.0 277.82 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  283.56 0.0 283.94 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  288.32 0.0 288.7 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 0.0 291.42 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 0.0 296.86 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  299.88 0.0 300.26 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 0.0 300.94 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.0 0.0 306.38 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.68 0.0 307.06 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 309.78 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  312.8 0.0 313.18 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.24 0.0 318.62 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  320.96 0.0 321.34 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  324.36 0.0 324.74 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 0.0 326.1 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 0.0 330.86 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.84 0.0 332.22 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  336.6 0.0 336.98 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  337.96 0.0 338.34 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 0.0 343.1 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  346.8 0.0 347.18 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  349.52 0.0 349.9 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.2 0.0 350.58 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  356.32 0.0 356.7 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.04 0.0 359.42 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  361.76 0.0 362.14 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.16 0.0 365.54 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.88 0.0 368.26 1.06 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  371.28 0.0 371.66 1.06 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  374.0 0.0 374.38 1.06 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  375.36 0.0 375.74 1.06 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  378.76 0.0 379.14 1.06 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  381.48 0.0 381.86 1.06 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  387.6 0.0 387.98 1.06 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  389.64 0.0 390.02 1.06 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 0.0 393.42 1.06 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  395.76 0.0 396.14 1.06 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  399.84 0.0 400.22 1.06 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  400.52 0.0 400.9 1.06 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.96 0.0 406.34 1.06 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  406.64 0.0 407.02 1.06 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.08 0.0 412.46 1.06 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 0.0 413.14 1.06 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  414.8 0.0 415.18 1.06 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  422.28 0.0 422.66 1.06 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  424.32 0.0 424.7 1.06 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  425.0 0.0 425.38 1.06 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  431.12 0.0 431.5 1.06 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  431.8 0.0 432.18 1.06 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  436.56 0.0 436.94 1.06 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  437.92 0.0 438.3 1.06 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.68 0.0 443.06 1.06 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  446.08 0.0 446.46 1.06 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  448.8 0.0 449.18 1.06 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  452.88 0.0 453.26 1.06 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  455.6 0.0 455.98 1.06 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  458.32 0.0 458.7 1.06 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  459.68 0.0 460.06 1.06 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  464.44 0.0 464.82 1.06 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  465.8 0.0 466.18 1.06 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  471.24 0.0 471.62 1.06 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  474.64 0.0 475.02 1.06 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  477.36 0.0 477.74 1.06 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  478.04 0.0 478.42 1.06 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  481.44 0.0 481.82 1.06 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  484.84 0.0 485.22 1.06 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  487.56 0.0 487.94 1.06 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  490.28 0.0 490.66 1.06 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  495.72 0.0 496.1 1.06 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  499.8 0.0 500.18 1.06 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  500.48 0.0 500.86 1.06 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.24 0.0 505.62 1.06 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  506.6 0.0 506.98 1.06 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  511.36 0.0 511.74 1.06 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  512.72 0.0 513.1 1.06 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  517.48 0.0 517.86 1.06 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  522.24 0.0 522.62 1.06 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  524.28 0.0 524.66 1.06 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  524.96 0.0 525.34 1.06 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.4 0.0 530.78 1.06 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  531.08 0.0 531.46 1.06 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  536.52 0.0 536.9 1.06 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  539.92 0.0 540.3 1.06 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  542.64 0.0 543.02 1.06 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  546.04 0.0 546.42 1.06 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  548.76 0.0 549.14 1.06 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  552.16 0.0 552.54 1.06 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  554.88 0.0 555.26 1.06 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  558.28 0.0 558.66 1.06 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  559.64 0.0 560.02 1.06 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  564.4 0.0 564.78 1.06 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  565.76 0.0 566.14 1.06 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  570.52 0.0 570.9 1.06 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  574.6 0.0 574.98 1.06 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  575.28 0.0 575.66 1.06 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  580.04 0.0 580.42 1.06 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  581.4 0.0 581.78 1.06 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  586.84 0.0 587.22 1.06 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  587.52 0.0 587.9 1.06 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  592.96 0.0 593.34 1.06 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  595.68 0.0 596.06 1.06 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  599.08 0.0 599.46 1.06 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  599.76 0.0 600.14 1.06 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  605.88 0.0 606.26 1.06 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  606.56 0.0 606.94 1.06 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.0 0.0 612.38 1.06 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 0.0 613.06 1.06 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  617.44 0.0 617.82 1.06 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  621.52 0.0 621.9 1.06 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  624.24 0.0 624.62 1.06 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  624.92 0.0 625.3 1.06 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  630.36 0.0 630.74 1.06 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  633.08 0.0 633.46 1.06 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  636.48 0.0 636.86 1.06 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  639.88 0.0 640.26 1.06 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  642.6 0.0 642.98 1.06 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  646.0 0.0 646.38 1.06 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  646.68 0.0 647.06 1.06 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  650.08 0.0 650.46 1.06 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  652.8 0.0 653.18 1.06 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  658.24 0.0 658.62 1.06 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  661.64 0.0 662.02 1.06 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  664.36 0.0 664.74 1.06 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  665.72 0.0 666.1 1.06 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  670.48 0.0 670.86 1.06 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  674.56 0.0 674.94 1.06 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  676.6 0.0 676.98 1.06 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  680.68 0.0 681.06 1.06 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  681.36 0.0 681.74 1.06 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  686.12 0.0 686.5 1.06 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  687.48 0.0 687.86 1.06 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  692.24 0.0 692.62 1.06 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  697.0 0.0 697.38 1.06 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  699.04 0.0 699.42 1.06 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  699.72 0.0 700.1 1.06 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  705.16 0.0 705.54 1.06 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  705.84 0.0 706.22 1.06 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  711.28 0.0 711.66 1.06 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  712.64 0.0 713.02 1.06 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  717.4 0.0 717.78 1.06 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  721.48 0.0 721.86 1.06 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  724.2 0.0 724.58 1.06 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  727.6 0.0 727.98 1.06 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  729.64 0.0 730.02 1.06 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  733.04 0.0 733.42 1.06 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  734.4 0.0 734.78 1.06 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  739.16 0.0 739.54 1.06 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  740.52 0.0 740.9 1.06 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  745.28 0.0 745.66 1.06 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  746.64 0.0 747.02 1.06 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  750.04 0.0 750.42 1.06 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  755.48 0.0 755.86 1.06 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  756.16 0.0 756.54 1.06 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  761.6 0.0 761.98 1.06 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  762.28 0.0 762.66 1.06 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  767.04 0.0 767.42 1.06 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  770.44 0.0 770.82 1.06 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  773.84 0.0 774.22 1.06 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  774.52 0.0 774.9 1.06 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  780.64 0.0 781.02 1.06 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  782.68 0.0 783.06 1.06 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  786.08 0.0 786.46 1.06 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  787.44 0.0 787.82 1.06 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  792.2 0.0 792.58 1.06 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  796.96 0.0 797.34 1.06 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  798.32 0.0 798.7 1.06 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  799.68 0.0 800.06 1.06 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  804.44 0.0 804.82 1.06 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  805.8 0.0 806.18 1.06 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  811.24 0.0 811.62 1.06 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  811.92 0.0 812.3 1.06 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  817.36 0.0 817.74 1.06 ;
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  820.76 0.0 821.14 1.06 ;
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  823.48 0.0 823.86 1.06 ;
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  826.88 0.0 827.26 1.06 ;
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  827.56 0.0 827.94 1.06 ;
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  830.96 0.0 831.34 1.06 ;
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  833.68 0.0 834.06 1.06 ;
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  839.12 0.0 839.5 1.06 ;
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  840.48 0.0 840.86 1.06 ;
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  845.24 0.0 845.62 1.06 ;
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  848.64 0.0 849.02 1.06 ;
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  851.36 0.0 851.74 1.06 ;
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  854.76 0.0 855.14 1.06 ;
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  856.12 0.0 856.5 1.06 ;
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  861.56 0.0 861.94 1.06 ;
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  862.24 0.0 862.62 1.06 ;
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  867.0 0.0 867.38 1.06 ;
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  870.4 0.0 870.78 1.06 ;
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  873.8 0.0 874.18 1.06 ;
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  874.48 0.0 874.86 1.06 ;
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  879.92 0.0 880.3 1.06 ;
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  880.6 0.0 880.98 1.06 ;
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  886.04 0.0 886.42 1.06 ;
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  886.72 0.0 887.1 1.06 ;
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  892.16 0.0 892.54 1.06 ;
      END
   END dout0[199]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 348.84 269.66 349.9 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 348.84 275.1 349.9 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 348.84 276.46 349.9 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 348.84 281.22 349.9 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  281.52 348.84 281.9 349.9 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  287.64 348.84 288.02 349.9 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 348.84 289.38 349.9 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  293.08 348.84 293.46 349.9 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  294.44 348.84 294.82 349.9 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  299.2 348.84 299.58 349.9 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 348.84 300.94 349.9 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.0 348.84 306.38 349.9 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.68 348.84 307.06 349.9 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 348.84 311.82 349.9 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  312.8 348.84 313.18 349.9 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 348.84 317.94 349.9 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  319.6 348.84 319.98 349.9 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  324.36 348.84 324.74 349.9 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 348.84 326.1 349.9 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 348.84 330.86 349.9 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.84 348.84 332.22 349.9 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  336.6 348.84 336.98 349.9 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  338.64 348.84 339.02 349.9 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 348.84 343.1 349.9 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  344.76 348.84 345.14 349.9 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  349.52 348.84 349.9 349.9 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.2 348.84 350.58 349.9 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  356.32 348.84 356.7 349.9 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  357.0 348.84 357.38 349.9 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  362.44 348.84 362.82 349.9 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  363.12 348.84 363.5 349.9 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  368.56 348.84 368.94 349.9 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  369.24 348.84 369.62 349.9 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  374.0 348.84 374.38 349.9 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  375.36 348.84 375.74 349.9 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  380.12 348.84 380.5 349.9 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  381.48 348.84 381.86 349.9 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  386.24 348.84 386.62 349.9 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  388.28 348.84 388.66 349.9 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 348.84 393.42 349.9 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  395.08 348.84 395.46 349.9 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  399.16 348.84 399.54 349.9 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  401.2 348.84 401.58 349.9 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.28 348.84 405.66 349.9 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  407.32 348.84 407.7 349.9 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.08 348.84 412.46 349.9 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 348.84 413.14 349.9 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 348.84 417.9 349.9 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  418.88 348.84 419.26 349.9 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  425.0 348.84 425.38 349.9 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  425.68 348.84 426.06 349.9 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  430.44 348.84 430.82 349.9 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  431.8 348.84 432.18 349.9 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  437.24 348.84 437.62 349.9 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  437.92 348.84 438.3 349.9 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  443.36 348.84 443.74 349.9 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  444.04 348.84 444.42 349.9 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  449.48 348.84 449.86 349.9 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  450.16 348.84 450.54 349.9 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 348.84 455.3 349.9 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  456.96 348.84 457.34 349.9 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  461.72 348.84 462.1 349.9 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  463.08 348.84 463.46 349.9 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  468.52 348.84 468.9 349.9 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  469.88 348.84 470.26 349.9 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  474.64 348.84 475.02 349.9 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  475.32 348.84 475.7 349.9 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  480.08 348.84 480.46 349.9 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  481.44 348.84 481.82 349.9 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  486.88 348.84 487.26 349.9 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  487.56 348.84 487.94 349.9 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 348.84 492.7 349.9 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  493.68 348.84 494.06 349.9 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  499.12 348.84 499.5 349.9 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  500.48 348.84 500.86 349.9 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.24 348.84 505.62 349.9 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  506.6 348.84 506.98 349.9 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  511.36 348.84 511.74 349.9 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  513.4 348.84 513.78 349.9 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  518.16 348.84 518.54 349.9 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  518.84 348.84 519.22 349.9 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  524.28 348.84 524.66 349.9 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  524.96 348.84 525.34 349.9 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.4 348.84 530.78 349.9 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  531.76 348.84 532.14 349.9 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  537.2 348.84 537.58 349.9 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  537.88 348.84 538.26 349.9 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  542.64 348.84 543.02 349.9 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  544.0 348.84 544.38 349.9 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  548.76 348.84 549.14 349.9 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  550.8 348.84 551.18 349.9 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  554.88 348.84 555.26 349.9 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  556.92 348.84 557.3 349.9 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  561.0 348.84 561.38 349.9 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  563.04 348.84 563.42 349.9 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  568.48 348.84 568.86 349.9 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  569.84 348.84 570.22 349.9 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  573.92 348.84 574.3 349.9 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  575.96 348.84 576.34 349.9 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  580.72 348.84 581.1 349.9 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  582.08 348.84 582.46 349.9 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  586.16 348.84 586.54 349.9 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  587.52 348.84 587.9 349.9 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  592.96 348.84 593.34 349.9 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  593.64 348.84 594.02 349.9 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  598.4 348.84 598.78 349.9 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  599.76 348.84 600.14 349.9 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  605.88 348.84 606.26 349.9 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  606.56 348.84 606.94 349.9 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  611.32 348.84 611.7 349.9 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 348.84 613.06 349.9 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  617.44 348.84 617.82 349.9 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  619.48 348.84 619.86 349.9 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  623.56 348.84 623.94 349.9 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  624.92 348.84 625.3 349.9 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  629.68 348.84 630.06 349.9 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  631.72 348.84 632.1 349.9 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  636.48 348.84 636.86 349.9 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  637.84 348.84 638.22 349.9 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  642.6 348.84 642.98 349.9 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  644.64 348.84 645.02 349.9 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  649.4 348.84 649.78 349.9 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  650.08 348.84 650.46 349.9 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  655.52 348.84 655.9 349.9 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  656.88 348.84 657.26 349.9 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  661.64 348.84 662.02 349.9 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  662.32 348.84 662.7 349.9 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  667.08 348.84 667.46 349.9 ;
      END
   END dout1[127]
   PIN dout1[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  668.44 348.84 668.82 349.9 ;
      END
   END dout1[128]
   PIN dout1[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  673.88 348.84 674.26 349.9 ;
      END
   END dout1[129]
   PIN dout1[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  675.92 348.84 676.3 349.9 ;
      END
   END dout1[130]
   PIN dout1[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  680.0 348.84 680.38 349.9 ;
      END
   END dout1[131]
   PIN dout1[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  682.04 348.84 682.42 349.9 ;
      END
   END dout1[132]
   PIN dout1[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  686.8 348.84 687.18 349.9 ;
      END
   END dout1[133]
   PIN dout1[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  688.16 348.84 688.54 349.9 ;
      END
   END dout1[134]
   PIN dout1[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  692.92 348.84 693.3 349.9 ;
      END
   END dout1[135]
   PIN dout1[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  693.6 348.84 693.98 349.9 ;
      END
   END dout1[136]
   PIN dout1[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  698.36 348.84 698.74 349.9 ;
      END
   END dout1[137]
   PIN dout1[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  699.72 348.84 700.1 349.9 ;
      END
   END dout1[138]
   PIN dout1[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  705.16 348.84 705.54 349.9 ;
      END
   END dout1[139]
   PIN dout1[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  705.84 348.84 706.22 349.9 ;
      END
   END dout1[140]
   PIN dout1[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  711.28 348.84 711.66 349.9 ;
      END
   END dout1[141]
   PIN dout1[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  712.64 348.84 713.02 349.9 ;
      END
   END dout1[142]
   PIN dout1[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  717.4 348.84 717.78 349.9 ;
      END
   END dout1[143]
   PIN dout1[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  718.76 348.84 719.14 349.9 ;
      END
   END dout1[144]
   PIN dout1[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  723.52 348.84 723.9 349.9 ;
      END
   END dout1[145]
   PIN dout1[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  725.56 348.84 725.94 349.9 ;
      END
   END dout1[146]
   PIN dout1[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  729.64 348.84 730.02 349.9 ;
      END
   END dout1[147]
   PIN dout1[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  731.68 348.84 732.06 349.9 ;
      END
   END dout1[148]
   PIN dout1[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  736.44 348.84 736.82 349.9 ;
      END
   END dout1[149]
   PIN dout1[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  737.12 348.84 737.5 349.9 ;
      END
   END dout1[150]
   PIN dout1[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  741.88 348.84 742.26 349.9 ;
      END
   END dout1[151]
   PIN dout1[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  744.6 348.84 744.98 349.9 ;
      END
   END dout1[152]
   PIN dout1[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  749.36 348.84 749.74 349.9 ;
      END
   END dout1[153]
   PIN dout1[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  750.72 348.84 751.1 349.9 ;
      END
   END dout1[154]
   PIN dout1[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  755.48 348.84 755.86 349.9 ;
      END
   END dout1[155]
   PIN dout1[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  756.16 348.84 756.54 349.9 ;
      END
   END dout1[156]
   PIN dout1[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  761.6 348.84 761.98 349.9 ;
      END
   END dout1[157]
   PIN dout1[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  762.28 348.84 762.66 349.9 ;
      END
   END dout1[158]
   PIN dout1[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  767.72 348.84 768.1 349.9 ;
      END
   END dout1[159]
   PIN dout1[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  768.4 348.84 768.78 349.9 ;
      END
   END dout1[160]
   PIN dout1[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  773.16 348.84 773.54 349.9 ;
      END
   END dout1[161]
   PIN dout1[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  774.52 348.84 774.9 349.9 ;
      END
   END dout1[162]
   PIN dout1[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  780.64 348.84 781.02 349.9 ;
      END
   END dout1[163]
   PIN dout1[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  781.32 348.84 781.7 349.9 ;
      END
   END dout1[164]
   PIN dout1[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  786.08 348.84 786.46 349.9 ;
      END
   END dout1[165]
   PIN dout1[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  788.12 348.84 788.5 349.9 ;
      END
   END dout1[166]
   PIN dout1[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  792.2 348.84 792.58 349.9 ;
      END
   END dout1[167]
   PIN dout1[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  793.56 348.84 793.94 349.9 ;
      END
   END dout1[168]
   PIN dout1[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  798.32 348.84 798.7 349.9 ;
      END
   END dout1[169]
   PIN dout1[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  800.36 348.84 800.74 349.9 ;
      END
   END dout1[170]
   PIN dout1[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  804.44 348.84 804.82 349.9 ;
      END
   END dout1[171]
   PIN dout1[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  806.48 348.84 806.86 349.9 ;
      END
   END dout1[172]
   PIN dout1[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  811.24 348.84 811.62 349.9 ;
      END
   END dout1[173]
   PIN dout1[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  811.92 348.84 812.3 349.9 ;
      END
   END dout1[174]
   PIN dout1[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  817.36 348.84 817.74 349.9 ;
      END
   END dout1[175]
   PIN dout1[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  819.4 348.84 819.78 349.9 ;
      END
   END dout1[176]
   PIN dout1[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  824.16 348.84 824.54 349.9 ;
      END
   END dout1[177]
   PIN dout1[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  824.84 348.84 825.22 349.9 ;
      END
   END dout1[178]
   PIN dout1[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  830.28 348.84 830.66 349.9 ;
      END
   END dout1[179]
   PIN dout1[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  830.96 348.84 831.34 349.9 ;
      END
   END dout1[180]
   PIN dout1[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  835.72 348.84 836.1 349.9 ;
      END
   END dout1[181]
   PIN dout1[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  837.08 348.84 837.46 349.9 ;
      END
   END dout1[182]
   PIN dout1[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  841.84 348.84 842.22 349.9 ;
      END
   END dout1[183]
   PIN dout1[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  843.2 348.84 843.58 349.9 ;
      END
   END dout1[184]
   PIN dout1[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  848.64 348.84 849.02 349.9 ;
      END
   END dout1[185]
   PIN dout1[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  850.0 348.84 850.38 349.9 ;
      END
   END dout1[186]
   PIN dout1[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  855.44 348.84 855.82 349.9 ;
      END
   END dout1[187]
   PIN dout1[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  856.12 348.84 856.5 349.9 ;
      END
   END dout1[188]
   PIN dout1[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  861.56 348.84 861.94 349.9 ;
      END
   END dout1[189]
   PIN dout1[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  862.92 348.84 863.3 349.9 ;
      END
   END dout1[190]
   PIN dout1[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  867.0 348.84 867.38 349.9 ;
      END
   END dout1[191]
   PIN dout1[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  869.04 348.84 869.42 349.9 ;
      END
   END dout1[192]
   PIN dout1[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  873.8 348.84 874.18 349.9 ;
      END
   END dout1[193]
   PIN dout1[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  874.48 348.84 874.86 349.9 ;
      END
   END dout1[194]
   PIN dout1[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  879.24 348.84 879.62 349.9 ;
      END
   END dout1[195]
   PIN dout1[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  880.6 348.84 880.98 349.9 ;
      END
   END dout1[196]
   PIN dout1[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  886.72 348.84 887.1 349.9 ;
      END
   END dout1[197]
   PIN dout1[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  887.4 348.84 887.78 349.9 ;
      END
   END dout1[198]
   PIN dout1[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  892.16 348.84 892.54 349.9 ;
      END
   END dout1[199]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1527.28 3.4 1529.02 346.5 ;
         LAYER met4 ;
         RECT  3.4 3.4 5.14 346.5 ;
         LAYER met3 ;
         RECT  3.4 344.76 1529.02 346.5 ;
         LAYER met3 ;
         RECT  3.4 3.4 1529.02 5.14 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 348.16 1532.42 349.9 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 349.9 ;
         LAYER met4 ;
         RECT  1530.68 0.0 1532.42 349.9 ;
         LAYER met3 ;
         RECT  0.0 0.0 1532.42 1.74 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 1531.8 349.28 ;
   LAYER  met2 ;
      RECT  0.62 0.62 1531.8 349.28 ;
   LAYER  met3 ;
      RECT  1.66 136.08 1531.8 137.66 ;
      RECT  0.62 139.02 1.66 144.92 ;
      RECT  1.66 137.66 2.8 344.16 ;
      RECT  1.66 344.16 2.8 347.1 ;
      RECT  2.8 137.66 1529.62 344.16 ;
      RECT  1529.62 137.66 1531.8 344.16 ;
      RECT  1529.62 344.16 1531.8 347.1 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 136.08 ;
      RECT  2.8 5.74 1529.62 136.08 ;
      RECT  1529.62 2.8 1531.8 5.74 ;
      RECT  1529.62 5.74 1531.8 136.08 ;
      RECT  0.62 146.5 1.66 347.56 ;
      RECT  1.66 347.1 2.8 347.56 ;
      RECT  2.8 347.1 1529.62 347.56 ;
      RECT  1529.62 347.1 1531.8 347.56 ;
      RECT  0.62 2.34 1.66 136.08 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 1529.62 2.8 ;
      RECT  1529.62 2.34 1531.8 2.8 ;
   LAYER  met4 ;
      RECT  352.32 1.66 353.9 349.28 ;
      RECT  383.14 0.62 386.32 1.66 ;
      RECT  895.86 0.62 900.4 1.66 ;
      RECT  901.98 0.62 906.52 1.66 ;
      RECT  908.1 0.62 911.96 1.66 ;
      RECT  913.54 0.62 918.08 1.66 ;
      RECT  919.66 0.62 923.52 1.66 ;
      RECT  925.1 0.62 930.32 1.66 ;
      RECT  931.9 0.62 936.44 1.66 ;
      RECT  938.02 0.62 941.2 1.66 ;
      RECT  942.78 0.62 947.32 1.66 ;
      RECT  948.9 0.62 952.76 1.66 ;
      RECT  954.34 0.62 958.88 1.66 ;
      RECT  960.46 0.62 965.0 1.66 ;
      RECT  972.02 0.62 977.24 1.66 ;
      RECT  978.82 0.62 982.0 1.66 ;
      RECT  983.58 0.62 988.8 1.66 ;
      RECT  990.38 0.62 994.24 1.66 ;
      RECT  995.82 0.62 1000.36 1.66 ;
      RECT  1001.94 0.62 1006.48 1.66 ;
      RECT  1008.06 0.62 1011.24 1.66 ;
      RECT  1012.82 0.62 1018.04 1.66 ;
      RECT  1019.62 0.62 1022.8 1.66 ;
      RECT  1024.38 0.62 1028.92 1.66 ;
      RECT  1030.5 0.62 1035.72 1.66 ;
      RECT  1037.3 0.62 1040.48 1.66 ;
      RECT  1042.06 0.62 1047.28 1.66 ;
      RECT  1048.86 0.62 1052.72 1.66 ;
      RECT  1054.3 0.62 1058.84 1.66 ;
      RECT  1060.42 0.62 1064.96 1.66 ;
      RECT  1066.54 0.62 1069.72 1.66 ;
      RECT  1071.3 0.62 1076.52 1.66 ;
      RECT  1078.1 0.62 1081.96 1.66 ;
      RECT  1083.54 0.62 1088.08 1.66 ;
      RECT  1089.66 0.62 1093.52 1.66 ;
      RECT  1095.1 0.62 1099.64 1.66 ;
      RECT  1101.22 0.62 1105.08 1.66 ;
      RECT  1106.66 0.62 1111.2 1.66 ;
      RECT  1112.78 0.62 1116.64 1.66 ;
      RECT  1118.22 0.62 1122.08 1.66 ;
      RECT  1123.66 0.62 1128.2 1.66 ;
      RECT  1129.78 0.62 1135.0 1.66 ;
      RECT  1136.58 0.62 1139.76 1.66 ;
      RECT  1141.34 0.62 1145.88 1.66 ;
      RECT  1147.46 0.62 1152.0 1.66 ;
      RECT  1153.58 0.62 1158.12 1.66 ;
      RECT  1159.7 0.62 1162.88 1.66 ;
      RECT  1164.46 0.62 1169.0 1.66 ;
      RECT  1170.58 0.62 1175.12 1.66 ;
      RECT  1176.7 0.62 1180.56 1.66 ;
      RECT  1182.14 0.62 1186.68 1.66 ;
      RECT  1188.26 0.62 1193.48 1.66 ;
      RECT  1195.06 0.62 1198.24 1.66 ;
      RECT  1199.82 0.62 1205.04 1.66 ;
      RECT  1206.62 0.62 1209.8 1.66 ;
      RECT  1211.38 0.62 1216.6 1.66 ;
      RECT  1218.18 0.62 1222.72 1.66 ;
      RECT  1224.3 0.62 1228.16 1.66 ;
      RECT  1229.74 0.62 1233.6 1.66 ;
      RECT  1235.18 0.62 1239.72 1.66 ;
      RECT  1241.3 0.62 1245.16 1.66 ;
      RECT  1246.74 0.62 1250.6 1.66 ;
      RECT  1252.18 0.62 1256.72 1.66 ;
      RECT  1258.3 0.62 1263.52 1.66 ;
      RECT  1265.1 0.62 1268.96 1.66 ;
      RECT  1270.54 0.62 1274.4 1.66 ;
      RECT  1275.98 0.62 1280.52 1.66 ;
      RECT  1282.1 0.62 1286.64 1.66 ;
      RECT  1288.22 0.62 1291.4 1.66 ;
      RECT  1292.98 0.62 1298.2 1.66 ;
      RECT  1299.78 0.62 1303.64 1.66 ;
      RECT  1305.22 0.62 1309.08 1.66 ;
      RECT  1310.66 0.62 1315.2 1.66 ;
      RECT  1316.78 0.62 1322.0 1.66 ;
      RECT  1323.58 0.62 1326.76 1.66 ;
      RECT  1328.34 0.62 1332.88 1.66 ;
      RECT  1334.46 0.62 1338.32 1.66 ;
      RECT  1339.9 0.62 1345.12 1.66 ;
      RECT  1346.7 0.62 1349.88 1.66 ;
      RECT  1351.46 0.62 1356.68 1.66 ;
      RECT  1358.26 0.62 1361.44 1.66 ;
      RECT  1363.02 0.62 1368.24 1.66 ;
      RECT  1369.82 0.62 1373.68 1.66 ;
      RECT  1375.26 0.62 1379.12 1.66 ;
      RECT  1380.7 0.62 1385.24 1.66 ;
      RECT  1386.82 0.62 1391.36 1.66 ;
      RECT  1392.94 0.62 1396.8 1.66 ;
      RECT  1398.38 0.62 1402.92 1.66 ;
      RECT  1404.5 0.62 1408.36 1.66 ;
      RECT  1409.94 0.62 1414.48 1.66 ;
      RECT  1416.06 0.62 1421.28 1.66 ;
      RECT  1422.86 0.62 1426.72 1.66 ;
      RECT  1428.3 0.62 1432.84 1.66 ;
      RECT  1434.42 0.62 1438.28 1.66 ;
      RECT  1439.86 0.62 1444.4 1.66 ;
      RECT  1445.98 0.62 1449.84 1.66 ;
      RECT  1451.42 0.62 1455.96 1.66 ;
      RECT  1457.54 0.62 1462.08 1.66 ;
      RECT  1463.66 0.62 1466.84 1.66 ;
      RECT  1468.42 0.62 1473.64 1.66 ;
      RECT  1475.22 0.62 1478.4 1.66 ;
      RECT  1479.98 0.62 1485.2 1.66 ;
      RECT  1486.78 0.62 1489.96 1.66 ;
      RECT  1491.54 0.62 1496.76 1.66 ;
      RECT  1498.34 0.62 1502.88 1.66 ;
      RECT  1504.46 0.62 1508.32 1.66 ;
      RECT  1509.9 0.62 1513.76 1.66 ;
      RECT  196.6 1.66 198.18 348.24 ;
      RECT  198.18 1.66 352.32 348.24 ;
      RECT  194.1 348.24 194.56 349.28 ;
      RECT  353.9 1.66 966.36 348.24 ;
      RECT  966.36 1.66 967.94 348.24 ;
      RECT  968.62 0.62 970.44 1.66 ;
      RECT  968.62 348.24 1129.56 349.28 ;
      RECT  1131.14 348.24 1147.24 349.28 ;
      RECT  207.7 0.62 211.56 1.66 ;
      RECT  213.14 0.62 217.0 1.66 ;
      RECT  218.58 0.62 223.12 1.66 ;
      RECT  224.7 0.62 229.92 1.66 ;
      RECT  231.5 0.62 235.36 1.66 ;
      RECT  236.94 0.62 240.8 1.66 ;
      RECT  242.38 0.62 246.92 1.66 ;
      RECT  248.5 0.62 253.04 1.66 ;
      RECT  254.62 0.62 258.48 1.66 ;
      RECT  260.06 0.62 263.92 1.66 ;
      RECT  265.5 0.62 267.32 1.66 ;
      RECT  268.9 0.62 270.72 1.66 ;
      RECT  272.3 0.62 273.44 1.66 ;
      RECT  275.02 0.62 275.48 1.66 ;
      RECT  279.78 0.62 281.6 1.66 ;
      RECT  285.9 0.62 287.04 1.66 ;
      RECT  289.3 0.62 290.44 1.66 ;
      RECT  292.02 0.62 293.16 1.66 ;
      RECT  294.74 0.62 295.88 1.66 ;
      RECT  297.46 0.62 298.6 1.66 ;
      RECT  301.54 0.62 304.72 1.66 ;
      RECT  307.66 0.62 308.8 1.66 ;
      RECT  310.38 0.62 311.52 1.66 ;
      RECT  313.78 0.62 316.28 1.66 ;
      RECT  319.22 0.62 320.36 1.66 ;
      RECT  321.94 0.62 323.08 1.66 ;
      RECT  326.7 0.62 328.52 1.66 ;
      RECT  332.82 0.62 333.96 1.66 ;
      RECT  335.54 0.62 336.0 1.66 ;
      RECT  338.94 0.62 340.08 1.66 ;
      RECT  341.66 0.62 342.12 1.66 ;
      RECT  343.7 0.62 345.52 1.66 ;
      RECT  347.78 0.62 348.92 1.66 ;
      RECT  351.18 0.62 352.32 1.66 ;
      RECT  353.9 0.62 355.72 1.66 ;
      RECT  357.3 0.62 357.76 1.66 ;
      RECT  360.02 0.62 361.16 1.66 ;
      RECT  362.74 0.62 363.88 1.66 ;
      RECT  366.14 0.62 367.28 1.66 ;
      RECT  368.86 0.62 370.0 1.66 ;
      RECT  372.26 0.62 373.4 1.66 ;
      RECT  377.02 0.62 378.16 1.66 ;
      RECT  379.74 0.62 380.88 1.66 ;
      RECT  388.58 0.62 389.04 1.66 ;
      RECT  390.62 0.62 392.44 1.66 ;
      RECT  394.7 0.62 395.16 1.66 ;
      RECT  396.74 0.62 398.56 1.66 ;
      RECT  401.5 0.62 404.0 1.66 ;
      RECT  407.62 0.62 410.8 1.66 ;
      RECT  413.74 0.62 414.2 1.66 ;
      RECT  417.14 0.62 421.68 1.66 ;
      RECT  425.98 0.62 428.48 1.66 ;
      RECT  430.06 0.62 430.52 1.66 ;
      RECT  432.78 0.62 433.92 1.66 ;
      RECT  435.5 0.62 435.96 1.66 ;
      RECT  438.9 0.62 439.36 1.66 ;
      RECT  440.94 0.62 442.08 1.66 ;
      RECT  443.66 0.62 444.8 1.66 ;
      RECT  447.06 0.62 448.2 1.66 ;
      RECT  449.78 0.62 451.6 1.66 ;
      RECT  453.86 0.62 455.0 1.66 ;
      RECT  456.58 0.62 457.04 1.66 ;
      RECT  460.66 0.62 463.16 1.66 ;
      RECT  466.78 0.62 467.92 1.66 ;
      RECT  469.5 0.62 470.64 1.66 ;
      RECT  472.22 0.62 474.04 1.66 ;
      RECT  476.3 0.62 476.76 1.66 ;
      RECT  479.02 0.62 480.16 1.66 ;
      RECT  482.42 0.62 484.24 1.66 ;
      RECT  485.82 0.62 486.28 1.66 ;
      RECT  488.54 0.62 489.68 1.66 ;
      RECT  491.26 0.62 491.72 1.66 ;
      RECT  493.3 0.62 495.12 1.66 ;
      RECT  496.7 0.62 497.16 1.66 ;
      RECT  498.74 0.62 499.2 1.66 ;
      RECT  501.46 0.62 503.28 1.66 ;
      RECT  507.58 0.62 510.08 1.66 ;
      RECT  513.7 0.62 514.84 1.66 ;
      RECT  516.42 0.62 516.88 1.66 ;
      RECT  518.46 0.62 520.96 1.66 ;
      RECT  523.22 0.62 523.68 1.66 ;
      RECT  525.94 0.62 527.08 1.66 ;
      RECT  528.66 0.62 529.8 1.66 ;
      RECT  532.06 0.62 532.52 1.66 ;
      RECT  534.1 0.62 535.92 1.66 ;
      RECT  537.5 0.62 538.64 1.66 ;
      RECT  540.9 0.62 542.04 1.66 ;
      RECT  543.62 0.62 544.08 1.66 ;
      RECT  547.02 0.62 548.16 1.66 ;
      RECT  549.74 0.62 550.2 1.66 ;
      RECT  553.14 0.62 554.28 1.66 ;
      RECT  557.22 0.62 557.68 1.66 ;
      RECT  560.62 0.62 561.76 1.66 ;
      RECT  563.34 0.62 563.8 1.66 ;
      RECT  566.74 0.62 568.56 1.66 ;
      RECT  571.5 0.62 573.32 1.66 ;
      RECT  576.26 0.62 579.44 1.66 ;
      RECT  582.38 0.62 584.88 1.66 ;
      RECT  588.5 0.62 591.68 1.66 ;
      RECT  593.94 0.62 595.08 1.66 ;
      RECT  596.66 0.62 597.12 1.66 ;
      RECT  600.74 0.62 603.24 1.66 ;
      RECT  604.82 0.62 605.28 1.66 ;
      RECT  607.54 0.62 608.68 1.66 ;
      RECT  610.26 0.62 611.4 1.66 ;
      RECT  613.66 0.62 614.8 1.66 ;
      RECT  616.38 0.62 616.84 1.66 ;
      RECT  618.42 0.62 620.24 1.66 ;
      RECT  622.5 0.62 623.64 1.66 ;
      RECT  625.9 0.62 626.36 1.66 ;
      RECT  627.94 0.62 629.76 1.66 ;
      RECT  631.34 0.62 631.8 1.66 ;
      RECT  634.06 0.62 635.88 1.66 ;
      RECT  637.46 0.62 638.6 1.66 ;
      RECT  640.86 0.62 642.0 1.66 ;
      RECT  644.94 0.62 645.4 1.66 ;
      RECT  647.66 0.62 649.48 1.66 ;
      RECT  651.74 0.62 652.2 1.66 ;
      RECT  653.78 0.62 655.6 1.66 ;
      RECT  657.18 0.62 657.64 1.66 ;
      RECT  659.22 0.62 661.04 1.66 ;
      RECT  663.3 0.62 663.76 1.66 ;
      RECT  666.7 0.62 667.84 1.66 ;
      RECT  669.42 0.62 669.88 1.66 ;
      RECT  671.46 0.62 673.28 1.66 ;
      RECT  675.54 0.62 676.0 1.66 ;
      RECT  677.58 0.62 679.4 1.66 ;
      RECT  682.34 0.62 684.16 1.66 ;
      RECT  688.46 0.62 690.96 1.66 ;
      RECT  693.22 0.62 695.72 1.66 ;
      RECT  697.98 0.62 698.44 1.66 ;
      RECT  700.7 0.62 701.84 1.66 ;
      RECT  703.42 0.62 704.56 1.66 ;
      RECT  706.82 0.62 708.64 1.66 ;
      RECT  710.22 0.62 710.68 1.66 ;
      RECT  714.98 0.62 716.8 1.66 ;
      RECT  718.38 0.62 720.2 1.66 ;
      RECT  722.46 0.62 723.6 1.66 ;
      RECT  725.18 0.62 726.32 1.66 ;
      RECT  728.58 0.62 729.04 1.66 ;
      RECT  730.62 0.62 731.76 1.66 ;
      RECT  735.38 0.62 737.88 1.66 ;
      RECT  741.5 0.62 742.64 1.66 ;
      RECT  744.22 0.62 744.68 1.66 ;
      RECT  747.62 0.62 748.76 1.66 ;
      RECT  751.02 0.62 754.2 1.66 ;
      RECT  757.14 0.62 760.32 1.66 ;
      RECT  763.26 0.62 765.76 1.66 ;
      RECT  768.02 0.62 769.84 1.66 ;
      RECT  771.42 0.62 771.88 1.66 ;
      RECT  775.5 0.62 778.0 1.66 ;
      RECT  779.58 0.62 780.04 1.66 ;
      RECT  781.62 0.62 782.08 1.66 ;
      RECT  785.02 0.62 785.48 1.66 ;
      RECT  788.42 0.62 789.56 1.66 ;
      RECT  791.14 0.62 791.6 1.66 ;
      RECT  793.18 0.62 795.68 1.66 ;
      RECT  800.66 0.62 801.8 1.66 ;
      RECT  803.38 0.62 803.84 1.66 ;
      RECT  806.78 0.62 807.92 1.66 ;
      RECT  809.5 0.62 810.64 1.66 ;
      RECT  812.9 0.62 813.36 1.66 ;
      RECT  814.94 0.62 816.76 1.66 ;
      RECT  818.34 0.62 819.48 1.66 ;
      RECT  821.74 0.62 822.88 1.66 ;
      RECT  824.46 0.62 824.92 1.66 ;
      RECT  828.54 0.62 830.36 1.66 ;
      RECT  832.62 0.62 833.08 1.66 ;
      RECT  834.66 0.62 836.48 1.66 ;
      RECT  838.06 0.62 838.52 1.66 ;
      RECT  841.46 0.62 841.92 1.66 ;
      RECT  843.5 0.62 844.64 1.66 ;
      RECT  846.22 0.62 848.04 1.66 ;
      RECT  850.3 0.62 850.76 1.66 ;
      RECT  852.34 0.62 853.48 1.66 ;
      RECT  857.1 0.62 860.28 1.66 ;
      RECT  863.22 0.62 865.04 1.66 ;
      RECT  867.98 0.62 869.8 1.66 ;
      RECT  871.38 0.62 871.84 1.66 ;
      RECT  875.46 0.62 877.96 1.66 ;
      RECT  881.58 0.62 883.4 1.66 ;
      RECT  884.98 0.62 885.44 1.66 ;
      RECT  887.7 0.62 888.84 1.66 ;
      RECT  890.42 0.62 891.56 1.66 ;
      RECT  893.14 0.62 894.28 1.66 ;
      RECT  198.18 348.24 268.68 349.28 ;
      RECT  270.26 348.24 274.12 349.28 ;
      RECT  277.06 348.24 280.24 349.28 ;
      RECT  282.5 348.24 287.04 349.28 ;
      RECT  289.98 348.24 292.48 349.28 ;
      RECT  295.42 348.24 298.6 349.28 ;
      RECT  301.54 348.24 305.4 349.28 ;
      RECT  307.66 348.24 310.84 349.28 ;
      RECT  313.78 348.24 316.96 349.28 ;
      RECT  318.54 348.24 319.0 349.28 ;
      RECT  320.58 348.24 323.76 349.28 ;
      RECT  326.7 348.24 329.88 349.28 ;
      RECT  332.82 348.24 336.0 349.28 ;
      RECT  337.58 348.24 338.04 349.28 ;
      RECT  339.62 348.24 342.12 349.28 ;
      RECT  343.7 348.24 344.16 349.28 ;
      RECT  345.74 348.24 348.92 349.28 ;
      RECT  351.18 348.24 352.32 349.28 ;
      RECT  353.9 348.24 355.72 349.28 ;
      RECT  357.98 348.24 361.84 349.28 ;
      RECT  364.1 348.24 367.96 349.28 ;
      RECT  370.22 348.24 373.4 349.28 ;
      RECT  376.34 348.24 379.52 349.28 ;
      RECT  382.46 348.24 385.64 349.28 ;
      RECT  387.22 348.24 387.68 349.28 ;
      RECT  389.26 348.24 392.44 349.28 ;
      RECT  394.02 348.24 394.48 349.28 ;
      RECT  396.06 348.24 398.56 349.28 ;
      RECT  400.14 348.24 400.6 349.28 ;
      RECT  402.18 348.24 404.68 349.28 ;
      RECT  406.26 348.24 406.72 349.28 ;
      RECT  408.3 348.24 411.48 349.28 ;
      RECT  413.74 348.24 416.92 349.28 ;
      RECT  419.86 348.24 424.4 349.28 ;
      RECT  426.66 348.24 429.84 349.28 ;
      RECT  432.78 348.24 436.64 349.28 ;
      RECT  438.9 348.24 442.76 349.28 ;
      RECT  445.02 348.24 448.88 349.28 ;
      RECT  451.14 348.24 454.32 349.28 ;
      RECT  455.9 348.24 456.36 349.28 ;
      RECT  457.94 348.24 461.12 349.28 ;
      RECT  464.06 348.24 467.92 349.28 ;
      RECT  470.86 348.24 474.04 349.28 ;
      RECT  476.3 348.24 479.48 349.28 ;
      RECT  482.42 348.24 486.28 349.28 ;
      RECT  488.54 348.24 491.72 349.28 ;
      RECT  494.66 348.24 498.52 349.28 ;
      RECT  501.46 348.24 504.64 349.28 ;
      RECT  507.58 348.24 510.76 349.28 ;
      RECT  512.34 348.24 512.8 349.28 ;
      RECT  514.38 348.24 517.56 349.28 ;
      RECT  519.82 348.24 523.68 349.28 ;
      RECT  525.94 348.24 529.8 349.28 ;
      RECT  532.74 348.24 536.6 349.28 ;
      RECT  538.86 348.24 542.04 349.28 ;
      RECT  544.98 348.24 548.16 349.28 ;
      RECT  549.74 348.24 550.2 349.28 ;
      RECT  551.78 348.24 554.28 349.28 ;
      RECT  555.86 348.24 556.32 349.28 ;
      RECT  557.9 348.24 560.4 349.28 ;
      RECT  561.98 348.24 562.44 349.28 ;
      RECT  564.02 348.24 567.88 349.28 ;
      RECT  570.82 348.24 573.32 349.28 ;
      RECT  574.9 348.24 575.36 349.28 ;
      RECT  576.94 348.24 580.12 349.28 ;
      RECT  583.06 348.24 585.56 349.28 ;
      RECT  588.5 348.24 592.36 349.28 ;
      RECT  594.62 348.24 597.8 349.28 ;
      RECT  600.74 348.24 605.28 349.28 ;
      RECT  607.54 348.24 610.72 349.28 ;
      RECT  613.66 348.24 616.84 349.28 ;
      RECT  618.42 348.24 618.88 349.28 ;
      RECT  620.46 348.24 622.96 349.28 ;
      RECT  625.9 348.24 629.08 349.28 ;
      RECT  630.66 348.24 631.12 349.28 ;
      RECT  632.7 348.24 635.88 349.28 ;
      RECT  638.82 348.24 642.0 349.28 ;
      RECT  643.58 348.24 644.04 349.28 ;
      RECT  645.62 348.24 648.8 349.28 ;
      RECT  651.06 348.24 654.92 349.28 ;
      RECT  657.86 348.24 661.04 349.28 ;
      RECT  663.3 348.24 666.48 349.28 ;
      RECT  669.42 348.24 673.28 349.28 ;
      RECT  674.86 348.24 675.32 349.28 ;
      RECT  676.9 348.24 679.4 349.28 ;
      RECT  680.98 348.24 681.44 349.28 ;
      RECT  683.02 348.24 686.2 349.28 ;
      RECT  689.14 348.24 692.32 349.28 ;
      RECT  694.58 348.24 697.76 349.28 ;
      RECT  700.7 348.24 704.56 349.28 ;
      RECT  706.82 348.24 710.68 349.28 ;
      RECT  713.62 348.24 716.8 349.28 ;
      RECT  719.74 348.24 722.92 349.28 ;
      RECT  724.5 348.24 724.96 349.28 ;
      RECT  726.54 348.24 729.04 349.28 ;
      RECT  730.62 348.24 731.08 349.28 ;
      RECT  732.66 348.24 735.84 349.28 ;
      RECT  738.1 348.24 741.28 349.28 ;
      RECT  742.86 348.24 744.0 349.28 ;
      RECT  745.58 348.24 748.76 349.28 ;
      RECT  751.7 348.24 754.88 349.28 ;
      RECT  757.14 348.24 761.0 349.28 ;
      RECT  763.26 348.24 767.12 349.28 ;
      RECT  769.38 348.24 772.56 349.28 ;
      RECT  775.5 348.24 780.04 349.28 ;
      RECT  782.3 348.24 785.48 349.28 ;
      RECT  787.06 348.24 787.52 349.28 ;
      RECT  789.1 348.24 791.6 349.28 ;
      RECT  794.54 348.24 797.72 349.28 ;
      RECT  799.3 348.24 799.76 349.28 ;
      RECT  801.34 348.24 803.84 349.28 ;
      RECT  805.42 348.24 805.88 349.28 ;
      RECT  807.46 348.24 810.64 349.28 ;
      RECT  812.9 348.24 816.76 349.28 ;
      RECT  818.34 348.24 818.8 349.28 ;
      RECT  820.38 348.24 823.56 349.28 ;
      RECT  825.82 348.24 829.68 349.28 ;
      RECT  831.94 348.24 835.12 349.28 ;
      RECT  838.06 348.24 841.24 349.28 ;
      RECT  844.18 348.24 848.04 349.28 ;
      RECT  850.98 348.24 854.84 349.28 ;
      RECT  857.1 348.24 860.96 349.28 ;
      RECT  863.9 348.24 866.4 349.28 ;
      RECT  867.98 348.24 868.44 349.28 ;
      RECT  870.02 348.24 873.2 349.28 ;
      RECT  875.46 348.24 878.64 349.28 ;
      RECT  881.58 348.24 886.12 349.28 ;
      RECT  888.38 348.24 891.56 349.28 ;
      RECT  893.14 348.24 965.68 349.28 ;
      RECT  967.94 1.66 1526.68 2.8 ;
      RECT  967.94 2.8 1526.68 347.1 ;
      RECT  967.94 347.1 1526.68 348.24 ;
      RECT  1526.68 1.66 1529.62 2.8 ;
      RECT  1526.68 347.1 1529.62 348.24 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 347.1 5.74 348.24 ;
      RECT  5.74 1.66 196.6 2.8 ;
      RECT  5.74 2.8 196.6 347.1 ;
      RECT  5.74 347.1 196.6 348.24 ;
      RECT  2.34 348.24 191.84 349.28 ;
      RECT  2.34 0.62 206.12 1.66 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 347.1 ;
      RECT  2.34 347.1 2.8 348.24 ;
      RECT  1515.34 0.62 1530.08 1.66 ;
      RECT  1148.82 348.24 1530.08 349.28 ;
      RECT  1529.62 1.66 1530.08 2.8 ;
      RECT  1529.62 2.8 1530.08 347.1 ;
      RECT  1529.62 347.1 1530.08 348.24 ;
   END
END    sky130_sram_1kbytes_1rw1r_200x48_8
END    LIBRARY
