VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_0kbytes_1rw1r_64x32_8
   CLASS BLOCK ;
   SIZE 535.54 BY 220.02 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  155.04 0.0 155.42 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 0.0 162.22 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 0.0 166.98 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 0.0 173.78 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 0.0 179.22 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  190.4 0.0 190.78 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.84 0.0 196.22 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 0.0 202.34 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.08 0.0 208.46 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  213.52 0.0 213.9 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  220.32 0.0 220.7 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  225.08 0.0 225.46 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  237.32 0.0 237.7 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  260.44 0.0 260.82 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 0.0 266.26 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 0.0 273.06 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 0.0 278.5 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.56 0.0 283.94 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.68 0.0 290.06 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.8 0.0 296.18 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 0.0 301.62 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  307.36 0.0 307.74 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  312.8 0.0 313.18 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  318.92 0.0 319.3 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  325.04 0.0 325.42 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  331.16 0.0 331.54 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  336.6 0.0 336.98 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 0.0 343.1 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  348.84 0.0 349.22 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  353.6 0.0 353.98 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  359.72 0.0 360.1 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  365.16 0.0 365.54 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 0.0 372.34 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 0.0 377.78 1.06 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  383.52 0.0 383.9 1.06 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  389.64 0.0 390.02 1.06 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  395.08 0.0 395.46 1.06 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  401.2 0.0 401.58 1.06 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  406.64 0.0 407.02 1.06 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 0.0 413.14 1.06 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  418.2 0.0 418.58 1.06 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  423.64 0.0 424.02 1.06 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 0.0 430.14 1.06 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  435.88 0.0 436.26 1.06 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  441.32 0.0 441.7 1.06 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  447.44 0.0 447.82 1.06 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  453.56 0.0 453.94 1.06 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  459.0 0.0 459.38 1.06 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  464.44 0.0 464.82 1.06 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  470.56 0.0 470.94 1.06 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  476.68 0.0 477.06 1.06 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  482.12 0.0 482.5 1.06 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  488.24 0.0 488.62 1.06 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  494.36 0.0 494.74 1.06 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  500.48 0.0 500.86 1.06 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  505.92 0.0 506.3 1.06 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  512.04 0.0 512.42 1.06 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  518.16 0.0 518.54 1.06 ;
      END
   END din0[63]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.84 218.96 94.22 220.02 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.16 218.96 93.54 220.02 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.76 218.96 90.14 220.02 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  92.48 218.96 92.86 220.02 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.8 218.96 92.18 220.02 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  534.48 94.52 535.54 94.9 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  439.28 0.0 439.66 1.06 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  444.04 0.0 444.42 1.06 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  439.96 0.0 440.34 1.06 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  443.36 0.0 443.74 1.06 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 38.76 1.06 39.14 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  518.16 218.96 518.54 220.02 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 46.92 1.06 47.3 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 38.08 1.06 38.46 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  501.16 218.96 501.54 220.02 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  103.36 0.0 103.74 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.8 0.0 109.18 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  114.92 0.0 115.3 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  120.36 0.0 120.74 1.06 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.8 0.0 126.18 1.06 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.92 0.0 132.3 1.06 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 0.0 138.42 1.06 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 1.06 ;
      END
   END wmask0[7]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 0.0 169.02 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  174.76 0.0 175.14 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 0.0 179.9 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 0.0 182.62 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.64 0.0 186.02 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  188.36 0.0 188.74 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.8 0.0 194.18 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 0.0 198.26 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 0.0 209.82 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 0.0 210.5 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 0.0 222.74 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 0.0 223.42 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 0.0 228.86 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.16 0.0 229.54 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.92 0.0 234.3 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 0.0 235.66 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 0.0 239.06 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 0.0 244.5 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  246.84 0.0 247.22 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  249.56 0.0 249.94 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 0.0 253.34 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 0.0 256.74 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 0.0 257.42 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.16 0.0 263.54 1.06 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  268.6 0.0 268.98 1.06 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 0.0 275.1 1.06 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 0.0 281.22 1.06 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 0.0 284.62 1.06 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  285.6 0.0 285.98 1.06 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 0.0 290.74 1.06 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  293.76 0.0 294.14 1.06 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 0.0 296.86 1.06 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 1.06 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 0.0 302.98 1.06 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.96 0.0 304.34 1.06 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 309.78 1.06 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 0.0 310.46 1.06 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  315.52 0.0 315.9 1.06 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  319.6 0.0 319.98 1.06 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  321.64 0.0 322.02 1.06 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 0.0 323.38 1.06 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.44 0.0 328.82 1.06 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.84 0.0 332.22 1.06 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.56 0.0 334.94 1.06 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  337.28 0.0 337.66 1.06 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  340.0 0.0 340.38 1.06 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  343.4 0.0 343.78 1.06 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  344.76 0.0 345.14 1.06 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  349.52 0.0 349.9 1.06 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.88 0.0 351.26 1.06 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  355.64 0.0 356.02 1.06 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  357.0 0.0 357.38 1.06 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  360.4 0.0 360.78 1.06 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.84 0.0 366.22 1.06 ;
      END
   END dout0[63]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 218.96 166.98 220.02 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  171.36 218.96 171.74 220.02 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 218.96 173.1 220.02 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.16 218.96 178.54 220.02 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 218.96 179.9 220.02 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.28 218.96 184.66 220.02 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 218.96 186.7 220.02 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.08 218.96 191.46 220.02 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 218.96 192.14 220.02 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 218.96 197.58 220.02 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 218.96 198.94 220.02 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  202.64 218.96 203.02 220.02 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 218.96 205.06 220.02 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 218.96 210.5 220.02 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 218.96 211.86 220.02 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 218.96 216.62 220.02 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 218.96 217.3 220.02 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 218.96 222.74 220.02 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 218.96 223.42 220.02 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 218.96 228.86 220.02 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 218.96 230.22 220.02 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.6 218.96 234.98 220.02 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 218.96 235.66 220.02 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.04 218.96 240.42 220.02 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.08 218.96 242.46 220.02 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 218.96 247.9 220.02 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 218.96 248.58 220.02 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 218.96 253.34 220.02 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 218.96 255.38 220.02 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.08 218.96 259.46 220.02 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 218.96 261.5 220.02 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.2 218.96 265.58 220.02 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.24 218.96 267.62 220.02 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  271.32 218.96 271.7 220.02 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 218.96 273.06 220.02 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  277.44 218.96 277.82 220.02 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  279.48 218.96 279.86 220.02 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 218.96 284.62 220.02 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 218.96 286.66 220.02 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 218.96 291.42 220.02 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.72 218.96 292.1 220.02 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 218.96 296.86 220.02 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 218.96 298.22 220.02 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 218.96 302.98 220.02 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.96 218.96 304.34 220.02 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 218.96 309.78 220.02 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 218.96 310.46 220.02 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  314.84 218.96 315.22 220.02 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 218.96 317.94 220.02 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  321.64 218.96 322.02 220.02 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 218.96 323.38 220.02 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  327.76 218.96 328.14 220.02 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.12 218.96 329.5 220.02 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  333.88 218.96 334.26 220.02 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.92 218.96 336.3 220.02 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  340.0 218.96 340.38 220.02 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.04 218.96 342.42 220.02 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  346.12 218.96 346.5 220.02 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  347.48 218.96 347.86 220.02 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  353.6 218.96 353.98 220.02 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 218.96 355.34 220.02 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.04 218.96 359.42 220.02 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  361.08 218.96 361.46 220.02 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.16 218.96 365.54 220.02 ;
      END
   END dout1[63]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.4 3.4 5.14 216.62 ;
         LAYER met3 ;
         RECT  3.4 214.88 532.14 216.62 ;
         LAYER met4 ;
         RECT  530.4 3.4 532.14 216.62 ;
         LAYER met3 ;
         RECT  3.4 3.4 532.14 5.14 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  533.8 0.0 535.54 220.02 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 220.02 ;
         LAYER met3 ;
         RECT  0.0 218.28 535.54 220.02 ;
         LAYER met3 ;
         RECT  0.0 0.0 535.54 1.74 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 534.92 219.4 ;
   LAYER  met2 ;
      RECT  0.62 0.62 534.92 219.4 ;
   LAYER  met3 ;
      RECT  0.62 93.92 533.88 95.5 ;
      RECT  1.66 38.16 533.88 39.74 ;
      RECT  1.66 39.74 533.88 93.92 ;
      RECT  0.62 39.74 1.66 46.32 ;
      RECT  0.62 47.9 1.66 93.92 ;
      RECT  0.62 95.5 2.8 214.28 ;
      RECT  0.62 214.28 2.8 217.22 ;
      RECT  2.8 95.5 532.74 214.28 ;
      RECT  532.74 95.5 533.88 214.28 ;
      RECT  532.74 214.28 533.88 217.22 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 38.16 ;
      RECT  2.8 5.74 532.74 38.16 ;
      RECT  532.74 2.8 533.88 5.74 ;
      RECT  532.74 5.74 533.88 38.16 ;
      RECT  533.88 95.5 534.92 217.68 ;
      RECT  0.62 217.22 2.8 217.68 ;
      RECT  2.8 217.22 532.74 217.68 ;
      RECT  532.74 217.22 533.88 217.68 ;
      RECT  533.88 2.34 534.92 93.92 ;
      RECT  0.62 2.34 1.66 37.48 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 532.74 2.8 ;
      RECT  532.74 2.34 533.88 2.8 ;
   LAYER  met4 ;
      RECT  149.68 1.66 151.26 219.4 ;
      RECT  151.26 0.62 154.44 1.66 ;
      RECT  156.02 0.62 161.24 1.66 ;
      RECT  162.82 0.62 166.0 1.66 ;
      RECT  372.94 0.62 376.8 1.66 ;
      RECT  378.38 0.62 382.92 1.66 ;
      RECT  384.5 0.62 389.04 1.66 ;
      RECT  390.62 0.62 394.48 1.66 ;
      RECT  396.06 0.62 400.6 1.66 ;
      RECT  402.18 0.62 406.04 1.66 ;
      RECT  407.62 0.62 412.16 1.66 ;
      RECT  413.74 0.62 417.6 1.66 ;
      RECT  419.18 0.62 423.04 1.66 ;
      RECT  424.62 0.62 429.16 1.66 ;
      RECT  430.74 0.62 435.28 1.66 ;
      RECT  448.42 0.62 452.96 1.66 ;
      RECT  454.54 0.62 458.4 1.66 ;
      RECT  459.98 0.62 463.84 1.66 ;
      RECT  465.42 0.62 469.96 1.66 ;
      RECT  471.54 0.62 476.08 1.66 ;
      RECT  477.66 0.62 481.52 1.66 ;
      RECT  483.1 0.62 487.64 1.66 ;
      RECT  489.22 0.62 493.76 1.66 ;
      RECT  495.34 0.62 499.88 1.66 ;
      RECT  501.46 0.62 505.32 1.66 ;
      RECT  506.9 0.62 511.44 1.66 ;
      RECT  513.02 0.62 517.56 1.66 ;
      RECT  93.24 1.66 94.82 218.36 ;
      RECT  94.82 1.66 149.68 218.36 ;
      RECT  94.82 218.36 149.68 219.4 ;
      RECT  90.74 218.36 91.2 219.4 ;
      RECT  436.86 0.62 438.68 1.66 ;
      RECT  445.02 0.62 446.84 1.66 ;
      RECT  442.3 0.62 442.76 1.66 ;
      RECT  151.26 1.66 517.56 218.36 ;
      RECT  517.56 1.66 519.14 218.36 ;
      RECT  502.14 218.36 517.56 219.4 ;
      RECT  104.34 0.62 108.2 1.66 ;
      RECT  109.78 0.62 114.32 1.66 ;
      RECT  115.9 0.62 119.76 1.66 ;
      RECT  121.34 0.62 125.2 1.66 ;
      RECT  126.78 0.62 131.32 1.66 ;
      RECT  132.9 0.62 137.44 1.66 ;
      RECT  139.02 0.62 142.88 1.66 ;
      RECT  144.46 0.62 149.68 1.66 ;
      RECT  167.58 0.62 168.04 1.66 ;
      RECT  169.62 0.62 172.12 1.66 ;
      RECT  177.1 0.62 178.24 1.66 ;
      RECT  180.5 0.62 181.64 1.66 ;
      RECT  183.22 0.62 184.36 1.66 ;
      RECT  186.62 0.62 187.76 1.66 ;
      RECT  189.34 0.62 189.8 1.66 ;
      RECT  191.38 0.62 193.2 1.66 ;
      RECT  194.78 0.62 195.24 1.66 ;
      RECT  198.86 0.62 201.36 1.66 ;
      RECT  204.98 0.62 207.48 1.66 ;
      RECT  211.1 0.62 212.92 1.66 ;
      RECT  214.5 0.62 214.96 1.66 ;
      RECT  216.54 0.62 219.04 1.66 ;
      RECT  221.3 0.62 221.76 1.66 ;
      RECT  224.02 0.62 224.48 1.66 ;
      RECT  226.06 0.62 227.88 1.66 ;
      RECT  230.14 0.62 231.28 1.66 ;
      RECT  232.86 0.62 233.32 1.66 ;
      RECT  236.26 0.62 236.72 1.66 ;
      RECT  239.66 0.62 242.84 1.66 ;
      RECT  245.1 0.62 246.24 1.66 ;
      RECT  247.82 0.62 248.28 1.66 ;
      RECT  250.54 0.62 252.36 1.66 ;
      RECT  253.94 0.62 254.4 1.66 ;
      RECT  258.02 0.62 259.84 1.66 ;
      RECT  261.42 0.62 261.88 1.66 ;
      RECT  264.14 0.62 265.28 1.66 ;
      RECT  266.86 0.62 268.0 1.66 ;
      RECT  269.58 0.62 271.4 1.66 ;
      RECT  273.66 0.62 274.12 1.66 ;
      RECT  275.7 0.62 277.52 1.66 ;
      RECT  279.78 0.62 280.24 1.66 ;
      RECT  281.82 0.62 282.96 1.66 ;
      RECT  286.58 0.62 289.08 1.66 ;
      RECT  291.34 0.62 293.16 1.66 ;
      RECT  294.74 0.62 295.2 1.66 ;
      RECT  298.82 0.62 300.64 1.66 ;
      RECT  304.94 0.62 306.76 1.66 ;
      RECT  308.34 0.62 308.8 1.66 ;
      RECT  311.06 0.62 312.2 1.66 ;
      RECT  313.78 0.62 314.92 1.66 ;
      RECT  316.5 0.62 318.32 1.66 ;
      RECT  320.58 0.62 321.04 1.66 ;
      RECT  323.98 0.62 324.44 1.66 ;
      RECT  326.02 0.62 327.84 1.66 ;
      RECT  329.42 0.62 330.56 1.66 ;
      RECT  332.82 0.62 333.96 1.66 ;
      RECT  335.54 0.62 336.0 1.66 ;
      RECT  338.26 0.62 339.4 1.66 ;
      RECT  340.98 0.62 342.12 1.66 ;
      RECT  345.74 0.62 348.24 1.66 ;
      RECT  351.86 0.62 353.0 1.66 ;
      RECT  354.58 0.62 355.04 1.66 ;
      RECT  357.98 0.62 359.12 1.66 ;
      RECT  361.38 0.62 364.56 1.66 ;
      RECT  366.82 0.62 371.36 1.66 ;
      RECT  151.26 218.36 166.0 219.4 ;
      RECT  167.58 218.36 170.76 219.4 ;
      RECT  173.7 218.36 177.56 219.4 ;
      RECT  180.5 218.36 183.68 219.4 ;
      RECT  185.26 218.36 185.72 219.4 ;
      RECT  187.3 218.36 190.48 219.4 ;
      RECT  192.74 218.36 196.6 219.4 ;
      RECT  199.54 218.36 202.04 219.4 ;
      RECT  203.62 218.36 204.08 219.4 ;
      RECT  205.66 218.36 209.52 219.4 ;
      RECT  212.46 218.36 215.64 219.4 ;
      RECT  217.9 218.36 221.76 219.4 ;
      RECT  224.02 218.36 227.88 219.4 ;
      RECT  230.82 218.36 234.0 219.4 ;
      RECT  236.26 218.36 239.44 219.4 ;
      RECT  241.02 218.36 241.48 219.4 ;
      RECT  243.06 218.36 246.92 219.4 ;
      RECT  249.18 218.36 252.36 219.4 ;
      RECT  253.94 218.36 254.4 219.4 ;
      RECT  255.98 218.36 258.48 219.4 ;
      RECT  260.06 218.36 260.52 219.4 ;
      RECT  262.1 218.36 264.6 219.4 ;
      RECT  266.18 218.36 266.64 219.4 ;
      RECT  268.22 218.36 270.72 219.4 ;
      RECT  273.66 218.36 276.84 219.4 ;
      RECT  278.42 218.36 278.88 219.4 ;
      RECT  280.46 218.36 283.64 219.4 ;
      RECT  285.22 218.36 285.68 219.4 ;
      RECT  287.26 218.36 290.44 219.4 ;
      RECT  292.7 218.36 295.88 219.4 ;
      RECT  298.82 218.36 302.0 219.4 ;
      RECT  304.94 218.36 308.8 219.4 ;
      RECT  311.06 218.36 314.24 219.4 ;
      RECT  315.82 218.36 316.96 219.4 ;
      RECT  318.54 218.36 321.04 219.4 ;
      RECT  323.98 218.36 327.16 219.4 ;
      RECT  330.1 218.36 333.28 219.4 ;
      RECT  334.86 218.36 335.32 219.4 ;
      RECT  336.9 218.36 339.4 219.4 ;
      RECT  340.98 218.36 341.44 219.4 ;
      RECT  343.02 218.36 345.52 219.4 ;
      RECT  348.46 218.36 353.0 219.4 ;
      RECT  355.94 218.36 358.44 219.4 ;
      RECT  360.02 218.36 360.48 219.4 ;
      RECT  362.06 218.36 364.56 219.4 ;
      RECT  366.14 218.36 500.56 219.4 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 217.22 5.74 218.36 ;
      RECT  5.74 1.66 93.24 2.8 ;
      RECT  5.74 2.8 93.24 217.22 ;
      RECT  5.74 217.22 93.24 218.36 ;
      RECT  519.14 1.66 529.8 2.8 ;
      RECT  519.14 2.8 529.8 217.22 ;
      RECT  519.14 217.22 529.8 218.36 ;
      RECT  529.8 1.66 532.74 2.8 ;
      RECT  529.8 217.22 532.74 218.36 ;
      RECT  519.14 0.62 533.2 1.66 ;
      RECT  519.14 218.36 533.2 219.4 ;
      RECT  532.74 1.66 533.2 2.8 ;
      RECT  532.74 2.8 533.2 217.22 ;
      RECT  532.74 217.22 533.2 218.36 ;
      RECT  2.34 218.36 89.16 219.4 ;
      RECT  2.34 0.62 102.76 1.66 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 217.22 ;
      RECT  2.34 217.22 2.8 218.36 ;
   END
END    sky130_sram_0kbytes_1rw1r_64x32_8
END    LIBRARY
