module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vssa2,
    vdda2,
    vssa1,
    vdda1,
    vssd2,
    vccd2,
    vssd1,
    vccd1,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vssa2;
 input vdda2;
 input vssa1;
 input vdda1;
 input vssd2;
 input vccd2;
 input vssd1;
 input vccd1;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \efabless_subsystem.UNCONNECTED102 ;
 wire \efabless_subsystem._000_ ;
 wire \efabless_subsystem._001_ ;
 wire \efabless_subsystem._002_ ;
 wire \efabless_subsystem._003_ ;
 wire \efabless_subsystem._004_ ;
 wire \efabless_subsystem._005_ ;
 wire \efabless_subsystem._006_ ;
 wire \efabless_subsystem._007_ ;
 wire \efabless_subsystem._008_ ;
 wire \efabless_subsystem._009_ ;
 wire \efabless_subsystem._010_ ;
 wire \efabless_subsystem._011_ ;
 wire \efabless_subsystem._012_ ;
 wire \efabless_subsystem._013_ ;
 wire \efabless_subsystem._014_ ;
 wire \efabless_subsystem._015_ ;
 wire \efabless_subsystem._016_ ;
 wire \efabless_subsystem._017_ ;
 wire \efabless_subsystem._018_ ;
 wire \efabless_subsystem._019_ ;
 wire \efabless_subsystem._020_ ;
 wire \efabless_subsystem._021_ ;
 wire \efabless_subsystem._022_ ;
 wire \efabless_subsystem._023_ ;
 wire \efabless_subsystem._024_ ;
 wire \efabless_subsystem._025_ ;
 wire \efabless_subsystem._026_ ;
 wire \efabless_subsystem._027_ ;
 wire \efabless_subsystem._028_ ;
 wire \efabless_subsystem._029_ ;
 wire \efabless_subsystem._030_ ;
 wire \efabless_subsystem._031_ ;
 wire \efabless_subsystem._032_ ;
 wire \efabless_subsystem._033_ ;
 wire \efabless_subsystem._034_ ;
 wire \efabless_subsystem._035_ ;
 wire \efabless_subsystem._036_ ;
 wire \efabless_subsystem._037_ ;
 wire \efabless_subsystem._038_ ;
 wire \efabless_subsystem._039_ ;
 wire \efabless_subsystem._040_ ;
 wire \efabless_subsystem._041_ ;
 wire \efabless_subsystem._042_ ;
 wire \efabless_subsystem._043_ ;
 wire \efabless_subsystem._044_ ;
 wire \efabless_subsystem._045_ ;
 wire \efabless_subsystem._046_ ;
 wire \efabless_subsystem._047_ ;
 wire \efabless_subsystem._048_ ;
 wire \efabless_subsystem._049_ ;
 wire \efabless_subsystem._050_ ;
 wire \efabless_subsystem._051_ ;
 wire \efabless_subsystem._052_ ;
 wire \efabless_subsystem._053_ ;
 wire \efabless_subsystem._054_ ;
 wire \efabless_subsystem._055_ ;
 wire \efabless_subsystem._056_ ;
 wire \efabless_subsystem._057_ ;
 wire \efabless_subsystem._058_ ;
 wire \efabless_subsystem._059_ ;
 wire \efabless_subsystem._060_ ;
 wire \efabless_subsystem._061_ ;
 wire \efabless_subsystem._062_ ;
 wire \efabless_subsystem._063_ ;
 wire \efabless_subsystem._064_ ;
 wire \efabless_subsystem._065_ ;
 wire \efabless_subsystem._066_ ;
 wire \efabless_subsystem._067_ ;
 wire \efabless_subsystem._068_ ;
 wire \efabless_subsystem._069_ ;
 wire \efabless_subsystem._070_ ;
 wire \efabless_subsystem._071_ ;
 wire \efabless_subsystem._072_ ;
 wire \efabless_subsystem._073_ ;
 wire \efabless_subsystem._074_ ;
 wire \efabless_subsystem._075_ ;
 wire \efabless_subsystem._076_ ;
 wire \efabless_subsystem._077_ ;
 wire \efabless_subsystem._078_ ;
 wire \efabless_subsystem._079_ ;
 wire \efabless_subsystem._080_ ;
 wire \efabless_subsystem._081_ ;
 wire \efabless_subsystem._082_ ;
 wire \efabless_subsystem._083_ ;
 wire \efabless_subsystem._084_ ;
 wire \efabless_subsystem._085_ ;
 wire \efabless_subsystem._086_ ;
 wire \efabless_subsystem._087_ ;
 wire \efabless_subsystem._088_ ;
 wire \efabless_subsystem._089_ ;
 wire \efabless_subsystem._090_ ;
 wire \efabless_subsystem._091_ ;
 wire \efabless_subsystem._092_ ;
 wire \efabless_subsystem._093_ ;
 wire \efabless_subsystem._094_ ;
 wire \efabless_subsystem._095_ ;
 wire \efabless_subsystem._096_ ;
 wire \efabless_subsystem._097_ ;
 wire \efabless_subsystem._098_ ;
 wire \efabless_subsystem._099_ ;
 wire \efabless_subsystem._100_ ;
 wire \efabless_subsystem._101_ ;
 wire \efabless_subsystem._102_ ;
 wire \efabless_subsystem._103_ ;
 wire \efabless_subsystem._104_ ;
 wire \efabless_subsystem._105_ ;
 wire \efabless_subsystem._106_ ;
 wire \efabless_subsystem._107_ ;
 wire \efabless_subsystem._108_ ;
 wire \efabless_subsystem._109_ ;
 wire \efabless_subsystem._110_ ;
 wire \efabless_subsystem._111_ ;
 wire \efabless_subsystem._112_ ;
 wire \efabless_subsystem._113_ ;
 wire \efabless_subsystem._114_ ;
 wire \efabless_subsystem._115_ ;
 wire \efabless_subsystem._116_ ;
 wire \efabless_subsystem._117_ ;
 wire \efabless_subsystem._118_ ;
 wire \efabless_subsystem._119_ ;
 wire \efabless_subsystem._120_ ;
 wire \efabless_subsystem._121_ ;
 wire \efabless_subsystem._122_ ;
 wire \efabless_subsystem._123_ ;
 wire \efabless_subsystem._124_ ;
 wire \efabless_subsystem._125_ ;
 wire \efabless_subsystem._126_ ;
 wire \efabless_subsystem._127_ ;
 wire \efabless_subsystem._128_ ;
 wire \efabless_subsystem._129_ ;
 wire \efabless_subsystem._130_ ;
 wire \efabless_subsystem._131_ ;
 wire \efabless_subsystem._132_ ;
 wire \efabless_subsystem._133_ ;
 wire \efabless_subsystem._134_ ;
 wire \efabless_subsystem._135_ ;
 wire \efabless_subsystem._136_ ;
 wire \efabless_subsystem._137_ ;
 wire \efabless_subsystem._138_ ;
 wire \efabless_subsystem._139_ ;
 wire \efabless_subsystem._140_ ;
 wire \efabless_subsystem._141_ ;
 wire \efabless_subsystem._142_ ;
 wire \efabless_subsystem._143_ ;
 wire \efabless_subsystem._144_ ;
 wire \efabless_subsystem._145_ ;
 wire \efabless_subsystem._146_ ;
 wire \efabless_subsystem._147_ ;
 wire \efabless_subsystem._148_ ;
 wire \efabless_subsystem._149_ ;
 wire \efabless_subsystem._150_ ;
 wire \efabless_subsystem._151_ ;
 wire \efabless_subsystem._152_ ;
 wire \efabless_subsystem._153_ ;
 wire \efabless_subsystem._154_ ;
 wire \efabless_subsystem._155_ ;
 wire \efabless_subsystem._156_ ;
 wire \efabless_subsystem._157_ ;
 wire \efabless_subsystem._158_ ;
 wire \efabless_subsystem._159_ ;
 wire \efabless_subsystem._160_ ;
 wire \efabless_subsystem._161_ ;
 wire \efabless_subsystem._162_ ;
 wire \efabless_subsystem._163_ ;
 wire \efabless_subsystem._164_ ;
 wire \efabless_subsystem._165_ ;
 wire \efabless_subsystem._166_ ;
 wire \efabless_subsystem._167_ ;
 wire \efabless_subsystem._168_ ;
 wire \efabless_subsystem._169_ ;
 wire \efabless_subsystem._170_ ;
 wire \efabless_subsystem._171_ ;
 wire \efabless_subsystem._172_ ;
 wire \efabless_subsystem._173_ ;
 wire \efabless_subsystem._174_ ;
 wire \efabless_subsystem._175_ ;
 wire \efabless_subsystem._176_ ;
 wire \efabless_subsystem._177_ ;
 wire \efabless_subsystem._178_ ;
 wire \efabless_subsystem._179_ ;
 wire \efabless_subsystem._180_ ;
 wire \efabless_subsystem._181_ ;
 wire \efabless_subsystem._182_ ;
 wire \efabless_subsystem._183_ ;
 wire \efabless_subsystem._184_ ;
 wire \efabless_subsystem._185_ ;
 wire \efabless_subsystem._186_ ;
 wire \efabless_subsystem._187_ ;
 wire \efabless_subsystem._188_ ;
 wire \efabless_subsystem._189_ ;
 wire \efabless_subsystem._190_ ;
 wire \efabless_subsystem._191_ ;
 wire \efabless_subsystem._192_ ;
 wire \efabless_subsystem._193_ ;
 wire \efabless_subsystem._194_ ;
 wire \efabless_subsystem._195_ ;
 wire \efabless_subsystem._196_ ;
 wire \efabless_subsystem._197_ ;
 wire \efabless_subsystem._198_ ;
 wire \efabless_subsystem._199_ ;
 wire \efabless_subsystem._200_ ;
 wire \efabless_subsystem._201_ ;
 wire \efabless_subsystem._202_ ;
 wire \efabless_subsystem._203_ ;
 wire \efabless_subsystem._204_ ;
 wire \efabless_subsystem._205_ ;
 wire \efabless_subsystem._206_ ;
 wire \efabless_subsystem._207_ ;
 wire \efabless_subsystem._208_ ;
 wire \efabless_subsystem._209_ ;
 wire \efabless_subsystem._210_ ;
 wire \efabless_subsystem._211_ ;
 wire \efabless_subsystem._212_ ;
 wire \efabless_subsystem._213_ ;
 wire \efabless_subsystem._214_ ;
 wire \efabless_subsystem._215_ ;
 wire \efabless_subsystem._216_ ;
 wire \efabless_subsystem._217_ ;
 wire \efabless_subsystem._218_ ;
 wire \efabless_subsystem._219_ ;
 wire \efabless_subsystem._220_ ;
 wire \efabless_subsystem._221_ ;
 wire \efabless_subsystem._222_ ;
 wire \efabless_subsystem._223_ ;
 wire \efabless_subsystem.cfg_address[10] ;
 wire \efabless_subsystem.cfg_address[11] ;
 wire \efabless_subsystem.cfg_address[12] ;
 wire \efabless_subsystem.cfg_address[13] ;
 wire \efabless_subsystem.cfg_address[14] ;
 wire \efabless_subsystem.cfg_address[15] ;
 wire \efabless_subsystem.cfg_address[16] ;
 wire \efabless_subsystem.cfg_address[17] ;
 wire \efabless_subsystem.cfg_address[18] ;
 wire \efabless_subsystem.cfg_address[19] ;
 wire \efabless_subsystem.cfg_address[20] ;
 wire \efabless_subsystem.cfg_address[21] ;
 wire \efabless_subsystem.cfg_address[22] ;
 wire \efabless_subsystem.cfg_address[23] ;
 wire \efabless_subsystem.cfg_address[2] ;
 wire \efabless_subsystem.cfg_address[3] ;
 wire \efabless_subsystem.cfg_address[4] ;
 wire \efabless_subsystem.cfg_address[5] ;
 wire \efabless_subsystem.cfg_address[6] ;
 wire \efabless_subsystem.cfg_address[7] ;
 wire \efabless_subsystem.cfg_address[8] ;
 wire \efabless_subsystem.cfg_address[9] ;
 wire \efabless_subsystem.cfg_data_in[0] ;
 wire \efabless_subsystem.cfg_data_in[10] ;
 wire \efabless_subsystem.cfg_data_in[11] ;
 wire \efabless_subsystem.cfg_data_in[12] ;
 wire \efabless_subsystem.cfg_data_in[13] ;
 wire \efabless_subsystem.cfg_data_in[14] ;
 wire \efabless_subsystem.cfg_data_in[15] ;
 wire \efabless_subsystem.cfg_data_in[16] ;
 wire \efabless_subsystem.cfg_data_in[17] ;
 wire \efabless_subsystem.cfg_data_in[18] ;
 wire \efabless_subsystem.cfg_data_in[19] ;
 wire \efabless_subsystem.cfg_data_in[1] ;
 wire \efabless_subsystem.cfg_data_in[20] ;
 wire \efabless_subsystem.cfg_data_in[21] ;
 wire \efabless_subsystem.cfg_data_in[22] ;
 wire \efabless_subsystem.cfg_data_in[23] ;
 wire \efabless_subsystem.cfg_data_in[24] ;
 wire \efabless_subsystem.cfg_data_in[25] ;
 wire \efabless_subsystem.cfg_data_in[26] ;
 wire \efabless_subsystem.cfg_data_in[27] ;
 wire \efabless_subsystem.cfg_data_in[28] ;
 wire \efabless_subsystem.cfg_data_in[29] ;
 wire \efabless_subsystem.cfg_data_in[2] ;
 wire \efabless_subsystem.cfg_data_in[30] ;
 wire \efabless_subsystem.cfg_data_in[31] ;
 wire \efabless_subsystem.cfg_data_in[3] ;
 wire \efabless_subsystem.cfg_data_in[4] ;
 wire \efabless_subsystem.cfg_data_in[5] ;
 wire \efabless_subsystem.cfg_data_in[6] ;
 wire \efabless_subsystem.cfg_data_in[7] ;
 wire \efabless_subsystem.cfg_data_in[8] ;
 wire \efabless_subsystem.cfg_data_in[9] ;
 wire \efabless_subsystem.cfg_done ;
 wire \efabless_subsystem.cfg_wmask[0] ;
 wire \efabless_subsystem.cfg_wmask[10] ;
 wire \efabless_subsystem.cfg_wmask[11] ;
 wire \efabless_subsystem.cfg_wmask[12] ;
 wire \efabless_subsystem.cfg_wmask[13] ;
 wire \efabless_subsystem.cfg_wmask[14] ;
 wire \efabless_subsystem.cfg_wmask[15] ;
 wire \efabless_subsystem.cfg_wmask[16] ;
 wire \efabless_subsystem.cfg_wmask[17] ;
 wire \efabless_subsystem.cfg_wmask[18] ;
 wire \efabless_subsystem.cfg_wmask[19] ;
 wire \efabless_subsystem.cfg_wmask[1] ;
 wire \efabless_subsystem.cfg_wmask[20] ;
 wire \efabless_subsystem.cfg_wmask[21] ;
 wire \efabless_subsystem.cfg_wmask[22] ;
 wire \efabless_subsystem.cfg_wmask[23] ;
 wire \efabless_subsystem.cfg_wmask[24] ;
 wire \efabless_subsystem.cfg_wmask[25] ;
 wire \efabless_subsystem.cfg_wmask[26] ;
 wire \efabless_subsystem.cfg_wmask[27] ;
 wire \efabless_subsystem.cfg_wmask[28] ;
 wire \efabless_subsystem.cfg_wmask[29] ;
 wire \efabless_subsystem.cfg_wmask[2] ;
 wire \efabless_subsystem.cfg_wmask[30] ;
 wire \efabless_subsystem.cfg_wmask[31] ;
 wire \efabless_subsystem.cfg_wmask[3] ;
 wire \efabless_subsystem.cfg_wmask[4] ;
 wire \efabless_subsystem.cfg_wmask[5] ;
 wire \efabless_subsystem.cfg_wmask[6] ;
 wire \efabless_subsystem.cfg_wmask[7] ;
 wire \efabless_subsystem.cfg_wmask[8] ;
 wire \efabless_subsystem.cfg_wmask[9] ;
 wire \efabless_subsystem.cfg_wren ;
 wire \efabless_subsystem.compute_controller_i._0000_ ;
 wire \efabless_subsystem.compute_controller_i._0001_ ;
 wire \efabless_subsystem.compute_controller_i._0002_ ;
 wire \efabless_subsystem.compute_controller_i._0003_ ;
 wire \efabless_subsystem.compute_controller_i._0004_ ;
 wire \efabless_subsystem.compute_controller_i._0005_ ;
 wire \efabless_subsystem.compute_controller_i._0006_ ;
 wire \efabless_subsystem.compute_controller_i._0007_ ;
 wire \efabless_subsystem.compute_controller_i._0008_ ;
 wire \efabless_subsystem.compute_controller_i._0009_ ;
 wire \efabless_subsystem.compute_controller_i._0010_ ;
 wire \efabless_subsystem.compute_controller_i._0011_ ;
 wire \efabless_subsystem.compute_controller_i._0012_ ;
 wire \efabless_subsystem.compute_controller_i._0013_ ;
 wire \efabless_subsystem.compute_controller_i._0014_ ;
 wire \efabless_subsystem.compute_controller_i._0015_ ;
 wire \efabless_subsystem.compute_controller_i._0016_ ;
 wire \efabless_subsystem.compute_controller_i._0017_ ;
 wire \efabless_subsystem.compute_controller_i._0018_ ;
 wire \efabless_subsystem.compute_controller_i._0019_ ;
 wire \efabless_subsystem.compute_controller_i._0020_ ;
 wire \efabless_subsystem.compute_controller_i._0021_ ;
 wire \efabless_subsystem.compute_controller_i._0022_ ;
 wire \efabless_subsystem.compute_controller_i._0023_ ;
 wire \efabless_subsystem.compute_controller_i._0024_ ;
 wire \efabless_subsystem.compute_controller_i._0025_ ;
 wire \efabless_subsystem.compute_controller_i._0026_ ;
 wire \efabless_subsystem.compute_controller_i._0027_ ;
 wire \efabless_subsystem.compute_controller_i._0028_ ;
 wire \efabless_subsystem.compute_controller_i._0029_ ;
 wire \efabless_subsystem.compute_controller_i._0030_ ;
 wire \efabless_subsystem.compute_controller_i._0031_ ;
 wire \efabless_subsystem.compute_controller_i._0032_ ;
 wire \efabless_subsystem.compute_controller_i._0033_ ;
 wire \efabless_subsystem.compute_controller_i._0034_ ;
 wire \efabless_subsystem.compute_controller_i._0035_ ;
 wire \efabless_subsystem.compute_controller_i._0036_ ;
 wire \efabless_subsystem.compute_controller_i._0037_ ;
 wire \efabless_subsystem.compute_controller_i._0038_ ;
 wire \efabless_subsystem.compute_controller_i._0039_ ;
 wire \efabless_subsystem.compute_controller_i._0040_ ;
 wire \efabless_subsystem.compute_controller_i._0041_ ;
 wire \efabless_subsystem.compute_controller_i._0042_ ;
 wire \efabless_subsystem.compute_controller_i._0043_ ;
 wire \efabless_subsystem.compute_controller_i._0044_ ;
 wire \efabless_subsystem.compute_controller_i._0045_ ;
 wire \efabless_subsystem.compute_controller_i._0046_ ;
 wire \efabless_subsystem.compute_controller_i._0047_ ;
 wire \efabless_subsystem.compute_controller_i._0048_ ;
 wire \efabless_subsystem.compute_controller_i._0049_ ;
 wire \efabless_subsystem.compute_controller_i._0050_ ;
 wire \efabless_subsystem.compute_controller_i._0051_ ;
 wire \efabless_subsystem.compute_controller_i._0052_ ;
 wire \efabless_subsystem.compute_controller_i._0053_ ;
 wire \efabless_subsystem.compute_controller_i._0054_ ;
 wire \efabless_subsystem.compute_controller_i._0055_ ;
 wire \efabless_subsystem.compute_controller_i._0056_ ;
 wire \efabless_subsystem.compute_controller_i._0057_ ;
 wire \efabless_subsystem.compute_controller_i._0058_ ;
 wire \efabless_subsystem.compute_controller_i._0059_ ;
 wire \efabless_subsystem.compute_controller_i._0060_ ;
 wire \efabless_subsystem.compute_controller_i._0061_ ;
 wire \efabless_subsystem.compute_controller_i._0062_ ;
 wire \efabless_subsystem.compute_controller_i._0063_ ;
 wire \efabless_subsystem.compute_controller_i._0064_ ;
 wire \efabless_subsystem.compute_controller_i._0065_ ;
 wire \efabless_subsystem.compute_controller_i._0066_ ;
 wire \efabless_subsystem.compute_controller_i._0067_ ;
 wire \efabless_subsystem.compute_controller_i._0068_ ;
 wire \efabless_subsystem.compute_controller_i._0069_ ;
 wire \efabless_subsystem.compute_controller_i._0070_ ;
 wire \efabless_subsystem.compute_controller_i._0071_ ;
 wire \efabless_subsystem.compute_controller_i._0072_ ;
 wire \efabless_subsystem.compute_controller_i._0073_ ;
 wire \efabless_subsystem.compute_controller_i._0074_ ;
 wire \efabless_subsystem.compute_controller_i._0075_ ;
 wire \efabless_subsystem.compute_controller_i._0076_ ;
 wire \efabless_subsystem.compute_controller_i._0077_ ;
 wire \efabless_subsystem.compute_controller_i._0078_ ;
 wire \efabless_subsystem.compute_controller_i._0079_ ;
 wire \efabless_subsystem.compute_controller_i._0080_ ;
 wire \efabless_subsystem.compute_controller_i._0081_ ;
 wire \efabless_subsystem.compute_controller_i._0082_ ;
 wire \efabless_subsystem.compute_controller_i._0083_ ;
 wire \efabless_subsystem.compute_controller_i._0084_ ;
 wire \efabless_subsystem.compute_controller_i._0085_ ;
 wire \efabless_subsystem.compute_controller_i._0086_ ;
 wire \efabless_subsystem.compute_controller_i._0087_ ;
 wire \efabless_subsystem.compute_controller_i._0088_ ;
 wire \efabless_subsystem.compute_controller_i._0089_ ;
 wire \efabless_subsystem.compute_controller_i._0090_ ;
 wire \efabless_subsystem.compute_controller_i._0091_ ;
 wire \efabless_subsystem.compute_controller_i._0092_ ;
 wire \efabless_subsystem.compute_controller_i._0093_ ;
 wire \efabless_subsystem.compute_controller_i._0094_ ;
 wire \efabless_subsystem.compute_controller_i._0095_ ;
 wire \efabless_subsystem.compute_controller_i._0096_ ;
 wire \efabless_subsystem.compute_controller_i._0097_ ;
 wire \efabless_subsystem.compute_controller_i._0098_ ;
 wire \efabless_subsystem.compute_controller_i._0099_ ;
 wire \efabless_subsystem.compute_controller_i._0100_ ;
 wire \efabless_subsystem.compute_controller_i._0101_ ;
 wire \efabless_subsystem.compute_controller_i._0102_ ;
 wire \efabless_subsystem.compute_controller_i._0103_ ;
 wire \efabless_subsystem.compute_controller_i._0104_ ;
 wire \efabless_subsystem.compute_controller_i._0105_ ;
 wire \efabless_subsystem.compute_controller_i._0106_ ;
 wire \efabless_subsystem.compute_controller_i._0108_ ;
 wire \efabless_subsystem.compute_controller_i._0110_ ;
 wire \efabless_subsystem.compute_controller_i._0111_ ;
 wire \efabless_subsystem.compute_controller_i._0113_ ;
 wire \efabless_subsystem.compute_controller_i._0114_ ;
 wire \efabless_subsystem.compute_controller_i._0116_ ;
 wire \efabless_subsystem.compute_controller_i._0118_ ;
 wire \efabless_subsystem.compute_controller_i._0120_ ;
 wire \efabless_subsystem.compute_controller_i._0123_ ;
 wire \efabless_subsystem.compute_controller_i._0124_ ;
 wire \efabless_subsystem.compute_controller_i._0126_ ;
 wire \efabless_subsystem.compute_controller_i._0128_ ;
 wire \efabless_subsystem.compute_controller_i._0129_ ;
 wire \efabless_subsystem.compute_controller_i._0130_ ;
 wire \efabless_subsystem.compute_controller_i._0131_ ;
 wire \efabless_subsystem.compute_controller_i._0132_ ;
 wire \efabless_subsystem.compute_controller_i._0133_ ;
 wire \efabless_subsystem.compute_controller_i._0134_ ;
 wire \efabless_subsystem.compute_controller_i._0135_ ;
 wire \efabless_subsystem.compute_controller_i._0136_ ;
 wire \efabless_subsystem.compute_controller_i._0137_ ;
 wire \efabless_subsystem.compute_controller_i._0138_ ;
 wire \efabless_subsystem.compute_controller_i._0139_ ;
 wire \efabless_subsystem.compute_controller_i._0140_ ;
 wire \efabless_subsystem.compute_controller_i._0141_ ;
 wire \efabless_subsystem.compute_controller_i._0142_ ;
 wire \efabless_subsystem.compute_controller_i._0143_ ;
 wire \efabless_subsystem.compute_controller_i._0144_ ;
 wire \efabless_subsystem.compute_controller_i._0145_ ;
 wire \efabless_subsystem.compute_controller_i._0146_ ;
 wire \efabless_subsystem.compute_controller_i._0147_ ;
 wire \efabless_subsystem.compute_controller_i._0148_ ;
 wire \efabless_subsystem.compute_controller_i._0149_ ;
 wire \efabless_subsystem.compute_controller_i._0150_ ;
 wire \efabless_subsystem.compute_controller_i._0151_ ;
 wire \efabless_subsystem.compute_controller_i._0152_ ;
 wire \efabless_subsystem.compute_controller_i._0153_ ;
 wire \efabless_subsystem.compute_controller_i._0154_ ;
 wire \efabless_subsystem.compute_controller_i._0155_ ;
 wire \efabless_subsystem.compute_controller_i._0156_ ;
 wire \efabless_subsystem.compute_controller_i._0157_ ;
 wire \efabless_subsystem.compute_controller_i._0158_ ;
 wire \efabless_subsystem.compute_controller_i._0159_ ;
 wire \efabless_subsystem.compute_controller_i._0160_ ;
 wire \efabless_subsystem.compute_controller_i._0161_ ;
 wire \efabless_subsystem.compute_controller_i._0162_ ;
 wire \efabless_subsystem.compute_controller_i._0163_ ;
 wire \efabless_subsystem.compute_controller_i._0164_ ;
 wire \efabless_subsystem.compute_controller_i._0165_ ;
 wire \efabless_subsystem.compute_controller_i._0166_ ;
 wire \efabless_subsystem.compute_controller_i._0167_ ;
 wire \efabless_subsystem.compute_controller_i._0168_ ;
 wire \efabless_subsystem.compute_controller_i._0169_ ;
 wire \efabless_subsystem.compute_controller_i._0170_ ;
 wire \efabless_subsystem.compute_controller_i._0171_ ;
 wire \efabless_subsystem.compute_controller_i._0172_ ;
 wire \efabless_subsystem.compute_controller_i._0173_ ;
 wire \efabless_subsystem.compute_controller_i._0174_ ;
 wire \efabless_subsystem.compute_controller_i._0175_ ;
 wire \efabless_subsystem.compute_controller_i._0176_ ;
 wire \efabless_subsystem.compute_controller_i._0177_ ;
 wire \efabless_subsystem.compute_controller_i._0178_ ;
 wire \efabless_subsystem.compute_controller_i._0179_ ;
 wire \efabless_subsystem.compute_controller_i._0180_ ;
 wire \efabless_subsystem.compute_controller_i._0181_ ;
 wire \efabless_subsystem.compute_controller_i._0182_ ;
 wire \efabless_subsystem.compute_controller_i._0183_ ;
 wire \efabless_subsystem.compute_controller_i._0184_ ;
 wire \efabless_subsystem.compute_controller_i._0185_ ;
 wire \efabless_subsystem.compute_controller_i._0186_ ;
 wire \efabless_subsystem.compute_controller_i._0187_ ;
 wire \efabless_subsystem.compute_controller_i._0188_ ;
 wire \efabless_subsystem.compute_controller_i._0189_ ;
 wire \efabless_subsystem.compute_controller_i._0190_ ;
 wire \efabless_subsystem.compute_controller_i._0191_ ;
 wire \efabless_subsystem.compute_controller_i._0192_ ;
 wire \efabless_subsystem.compute_controller_i._0193_ ;
 wire \efabless_subsystem.compute_controller_i._0194_ ;
 wire \efabless_subsystem.compute_controller_i._0195_ ;
 wire \efabless_subsystem.compute_controller_i._0196_ ;
 wire \efabless_subsystem.compute_controller_i._0197_ ;
 wire \efabless_subsystem.compute_controller_i._0198_ ;
 wire \efabless_subsystem.compute_controller_i._0199_ ;
 wire \efabless_subsystem.compute_controller_i._0200_ ;
 wire \efabless_subsystem.compute_controller_i._0201_ ;
 wire \efabless_subsystem.compute_controller_i._0202_ ;
 wire \efabless_subsystem.compute_controller_i._0203_ ;
 wire \efabless_subsystem.compute_controller_i._0204_ ;
 wire \efabless_subsystem.compute_controller_i._0205_ ;
 wire \efabless_subsystem.compute_controller_i._0206_ ;
 wire \efabless_subsystem.compute_controller_i._0207_ ;
 wire \efabless_subsystem.compute_controller_i._0208_ ;
 wire \efabless_subsystem.compute_controller_i._0209_ ;
 wire \efabless_subsystem.compute_controller_i._0210_ ;
 wire \efabless_subsystem.compute_controller_i._0211_ ;
 wire \efabless_subsystem.compute_controller_i._0212_ ;
 wire \efabless_subsystem.compute_controller_i._0213_ ;
 wire \efabless_subsystem.compute_controller_i._0214_ ;
 wire \efabless_subsystem.compute_controller_i._0215_ ;
 wire \efabless_subsystem.compute_controller_i._0216_ ;
 wire \efabless_subsystem.compute_controller_i._0217_ ;
 wire \efabless_subsystem.compute_controller_i._0218_ ;
 wire \efabless_subsystem.compute_controller_i._0219_ ;
 wire \efabless_subsystem.compute_controller_i._0220_ ;
 wire \efabless_subsystem.compute_controller_i._0221_ ;
 wire \efabless_subsystem.compute_controller_i._0222_ ;
 wire \efabless_subsystem.compute_controller_i._0223_ ;
 wire \efabless_subsystem.compute_controller_i._0224_ ;
 wire \efabless_subsystem.compute_controller_i._0225_ ;
 wire \efabless_subsystem.compute_controller_i._0226_ ;
 wire \efabless_subsystem.compute_controller_i._0227_ ;
 wire \efabless_subsystem.compute_controller_i._0228_ ;
 wire \efabless_subsystem.compute_controller_i._0229_ ;
 wire \efabless_subsystem.compute_controller_i._0230_ ;
 wire \efabless_subsystem.compute_controller_i._0231_ ;
 wire \efabless_subsystem.compute_controller_i._0232_ ;
 wire \efabless_subsystem.compute_controller_i._0233_ ;
 wire \efabless_subsystem.compute_controller_i._0234_ ;
 wire \efabless_subsystem.compute_controller_i._0235_ ;
 wire \efabless_subsystem.compute_controller_i._0236_ ;
 wire \efabless_subsystem.compute_controller_i._0237_ ;
 wire \efabless_subsystem.compute_controller_i._0238_ ;
 wire \efabless_subsystem.compute_controller_i._0239_ ;
 wire \efabless_subsystem.compute_controller_i._0240_ ;
 wire \efabless_subsystem.compute_controller_i._0241_ ;
 wire \efabless_subsystem.compute_controller_i._0242_ ;
 wire \efabless_subsystem.compute_controller_i._0243_ ;
 wire \efabless_subsystem.compute_controller_i._0244_ ;
 wire \efabless_subsystem.compute_controller_i._0245_ ;
 wire \efabless_subsystem.compute_controller_i._0246_ ;
 wire \efabless_subsystem.compute_controller_i._0247_ ;
 wire \efabless_subsystem.compute_controller_i._0248_ ;
 wire \efabless_subsystem.compute_controller_i._0249_ ;
 wire \efabless_subsystem.compute_controller_i._0250_ ;
 wire \efabless_subsystem.compute_controller_i._0251_ ;
 wire \efabless_subsystem.compute_controller_i._0252_ ;
 wire \efabless_subsystem.compute_controller_i._0253_ ;
 wire \efabless_subsystem.compute_controller_i._0254_ ;
 wire \efabless_subsystem.compute_controller_i._0255_ ;
 wire \efabless_subsystem.compute_controller_i._0256_ ;
 wire \efabless_subsystem.compute_controller_i._0257_ ;
 wire \efabless_subsystem.compute_controller_i._0258_ ;
 wire \efabless_subsystem.compute_controller_i._0259_ ;
 wire \efabless_subsystem.compute_controller_i._0260_ ;
 wire \efabless_subsystem.compute_controller_i._0261_ ;
 wire \efabless_subsystem.compute_controller_i._0262_ ;
 wire \efabless_subsystem.compute_controller_i._0263_ ;
 wire \efabless_subsystem.compute_controller_i._0264_ ;
 wire \efabless_subsystem.compute_controller_i._0265_ ;
 wire \efabless_subsystem.compute_controller_i._0266_ ;
 wire \efabless_subsystem.compute_controller_i._0267_ ;
 wire \efabless_subsystem.compute_controller_i._0268_ ;
 wire \efabless_subsystem.compute_controller_i._0269_ ;
 wire \efabless_subsystem.compute_controller_i._0270_ ;
 wire \efabless_subsystem.compute_controller_i._0271_ ;
 wire \efabless_subsystem.compute_controller_i._0272_ ;
 wire \efabless_subsystem.compute_controller_i._0273_ ;
 wire \efabless_subsystem.compute_controller_i._0274_ ;
 wire \efabless_subsystem.compute_controller_i._0275_ ;
 wire \efabless_subsystem.compute_controller_i._0276_ ;
 wire \efabless_subsystem.compute_controller_i._0277_ ;
 wire \efabless_subsystem.compute_controller_i._0278_ ;
 wire \efabless_subsystem.compute_controller_i._0279_ ;
 wire \efabless_subsystem.compute_controller_i._0280_ ;
 wire \efabless_subsystem.compute_controller_i._0281_ ;
 wire \efabless_subsystem.compute_controller_i._0282_ ;
 wire \efabless_subsystem.compute_controller_i._0283_ ;
 wire \efabless_subsystem.compute_controller_i._0284_ ;
 wire \efabless_subsystem.compute_controller_i._0285_ ;
 wire \efabless_subsystem.compute_controller_i._0286_ ;
 wire \efabless_subsystem.compute_controller_i._0287_ ;
 wire \efabless_subsystem.compute_controller_i._0288_ ;
 wire \efabless_subsystem.compute_controller_i._0289_ ;
 wire \efabless_subsystem.compute_controller_i._0290_ ;
 wire \efabless_subsystem.compute_controller_i._0291_ ;
 wire \efabless_subsystem.compute_controller_i._0292_ ;
 wire \efabless_subsystem.compute_controller_i._0293_ ;
 wire \efabless_subsystem.compute_controller_i._0294_ ;
 wire \efabless_subsystem.compute_controller_i._0295_ ;
 wire \efabless_subsystem.compute_controller_i._0296_ ;
 wire \efabless_subsystem.compute_controller_i._0297_ ;
 wire \efabless_subsystem.compute_controller_i._0298_ ;
 wire \efabless_subsystem.compute_controller_i._0299_ ;
 wire \efabless_subsystem.compute_controller_i._0300_ ;
 wire \efabless_subsystem.compute_controller_i._0301_ ;
 wire \efabless_subsystem.compute_controller_i._0302_ ;
 wire \efabless_subsystem.compute_controller_i._0303_ ;
 wire \efabless_subsystem.compute_controller_i._0304_ ;
 wire \efabless_subsystem.compute_controller_i._0305_ ;
 wire \efabless_subsystem.compute_controller_i._0306_ ;
 wire \efabless_subsystem.compute_controller_i._0307_ ;
 wire \efabless_subsystem.compute_controller_i._0308_ ;
 wire \efabless_subsystem.compute_controller_i._0309_ ;
 wire \efabless_subsystem.compute_controller_i._0310_ ;
 wire \efabless_subsystem.compute_controller_i._0311_ ;
 wire \efabless_subsystem.compute_controller_i._0312_ ;
 wire \efabless_subsystem.compute_controller_i._0313_ ;
 wire \efabless_subsystem.compute_controller_i._0314_ ;
 wire \efabless_subsystem.compute_controller_i._0315_ ;
 wire \efabless_subsystem.compute_controller_i._0316_ ;
 wire \efabless_subsystem.compute_controller_i._0317_ ;
 wire \efabless_subsystem.compute_controller_i._0318_ ;
 wire \efabless_subsystem.compute_controller_i._0319_ ;
 wire \efabless_subsystem.compute_controller_i._0320_ ;
 wire \efabless_subsystem.compute_controller_i._0321_ ;
 wire \efabless_subsystem.compute_controller_i._0322_ ;
 wire \efabless_subsystem.compute_controller_i._0323_ ;
 wire \efabless_subsystem.compute_controller_i._0324_ ;
 wire \efabless_subsystem.compute_controller_i._0325_ ;
 wire \efabless_subsystem.compute_controller_i._0326_ ;
 wire \efabless_subsystem.compute_controller_i._0327_ ;
 wire \efabless_subsystem.compute_controller_i._0328_ ;
 wire \efabless_subsystem.compute_controller_i._0329_ ;
 wire \efabless_subsystem.compute_controller_i._0330_ ;
 wire \efabless_subsystem.compute_controller_i._0331_ ;
 wire \efabless_subsystem.compute_controller_i._0332_ ;
 wire \efabless_subsystem.compute_controller_i._0333_ ;
 wire \efabless_subsystem.compute_controller_i._0334_ ;
 wire \efabless_subsystem.compute_controller_i._0335_ ;
 wire \efabless_subsystem.compute_controller_i._0336_ ;
 wire \efabless_subsystem.compute_controller_i._0337_ ;
 wire \efabless_subsystem.compute_controller_i._0338_ ;
 wire \efabless_subsystem.compute_controller_i._0339_ ;
 wire \efabless_subsystem.compute_controller_i._0340_ ;
 wire \efabless_subsystem.compute_controller_i._0341_ ;
 wire \efabless_subsystem.compute_controller_i._0342_ ;
 wire \efabless_subsystem.compute_controller_i._0343_ ;
 wire \efabless_subsystem.compute_controller_i._0344_ ;
 wire \efabless_subsystem.compute_controller_i._0345_ ;
 wire \efabless_subsystem.compute_controller_i._0346_ ;
 wire \efabless_subsystem.compute_controller_i._0347_ ;
 wire \efabless_subsystem.compute_controller_i._0348_ ;
 wire \efabless_subsystem.compute_controller_i._0349_ ;
 wire \efabless_subsystem.compute_controller_i._0350_ ;
 wire \efabless_subsystem.compute_controller_i._0351_ ;
 wire \efabless_subsystem.compute_controller_i._0352_ ;
 wire \efabless_subsystem.compute_controller_i._0353_ ;
 wire \efabless_subsystem.compute_controller_i._0354_ ;
 wire \efabless_subsystem.compute_controller_i._0355_ ;
 wire \efabless_subsystem.compute_controller_i._0356_ ;
 wire \efabless_subsystem.compute_controller_i._0357_ ;
 wire \efabless_subsystem.compute_controller_i._0358_ ;
 wire \efabless_subsystem.compute_controller_i._0359_ ;
 wire \efabless_subsystem.compute_controller_i._0360_ ;
 wire \efabless_subsystem.compute_controller_i._0361_ ;
 wire \efabless_subsystem.compute_controller_i._0362_ ;
 wire \efabless_subsystem.compute_controller_i._0363_ ;
 wire \efabless_subsystem.compute_controller_i._0364_ ;
 wire \efabless_subsystem.compute_controller_i._0365_ ;
 wire \efabless_subsystem.compute_controller_i._0366_ ;
 wire \efabless_subsystem.compute_controller_i._0367_ ;
 wire \efabless_subsystem.compute_controller_i._0368_ ;
 wire \efabless_subsystem.compute_controller_i._0369_ ;
 wire \efabless_subsystem.compute_controller_i._0371_ ;
 wire \efabless_subsystem.compute_controller_i._0372_ ;
 wire \efabless_subsystem.compute_controller_i._0373_ ;
 wire \efabless_subsystem.compute_controller_i._0374_ ;
 wire \efabless_subsystem.compute_controller_i._0375_ ;
 wire \efabless_subsystem.compute_controller_i._0376_ ;
 wire \efabless_subsystem.compute_controller_i._0377_ ;
 wire \efabless_subsystem.compute_controller_i._0378_ ;
 wire \efabless_subsystem.compute_controller_i._0379_ ;
 wire \efabless_subsystem.compute_controller_i._0380_ ;
 wire \efabless_subsystem.compute_controller_i._0381_ ;
 wire \efabless_subsystem.compute_controller_i._0382_ ;
 wire \efabless_subsystem.compute_controller_i._0383_ ;
 wire \efabless_subsystem.compute_controller_i._0384_ ;
 wire \efabless_subsystem.compute_controller_i._0385_ ;
 wire \efabless_subsystem.compute_controller_i._0386_ ;
 wire \efabless_subsystem.compute_controller_i._0387_ ;
 wire \efabless_subsystem.compute_controller_i._0388_ ;
 wire \efabless_subsystem.compute_controller_i._0389_ ;
 wire \efabless_subsystem.compute_controller_i._0390_ ;
 wire \efabless_subsystem.compute_controller_i._0391_ ;
 wire \efabless_subsystem.compute_controller_i._0392_ ;
 wire \efabless_subsystem.compute_controller_i._0393_ ;
 wire \efabless_subsystem.compute_controller_i._0394_ ;
 wire \efabless_subsystem.compute_controller_i._0395_ ;
 wire \efabless_subsystem.compute_controller_i._0396_ ;
 wire \efabless_subsystem.compute_controller_i._0397_ ;
 wire \efabless_subsystem.compute_controller_i._0401_ ;
 wire \efabless_subsystem.compute_controller_i._0402_ ;
 wire \efabless_subsystem.compute_controller_i._0403_ ;
 wire \efabless_subsystem.compute_controller_i._0407_ ;
 wire \efabless_subsystem.compute_controller_i._0408_ ;
 wire \efabless_subsystem.compute_controller_i._0412_ ;
 wire \efabless_subsystem.compute_controller_i._0413_ ;
 wire \efabless_subsystem.compute_controller_i._0414_ ;
 wire \efabless_subsystem.compute_controller_i._0418_ ;
 wire \efabless_subsystem.compute_controller_i._0419_ ;
 wire \efabless_subsystem.compute_controller_i._0420_ ;
 wire \efabless_subsystem.compute_controller_i._0423_ ;
 wire \efabless_subsystem.compute_controller_i._0424_ ;
 wire \efabless_subsystem.compute_controller_i._0427_ ;
 wire \efabless_subsystem.compute_controller_i._0430_ ;
 wire \efabless_subsystem.compute_controller_i._0431_ ;
 wire \efabless_subsystem.compute_controller_i._0435_ ;
 wire \efabless_subsystem.compute_controller_i._0436_ ;
 wire \efabless_subsystem.compute_controller_i._0439_ ;
 wire \efabless_subsystem.compute_controller_i._0440_ ;
 wire \efabless_subsystem.compute_controller_i._0443_ ;
 wire \efabless_subsystem.compute_controller_i._0444_ ;
 wire \efabless_subsystem.compute_controller_i._0447_ ;
 wire \efabless_subsystem.compute_controller_i._0448_ ;
 wire \efabless_subsystem.compute_controller_i._0450_ ;
 wire \efabless_subsystem.compute_controller_i._0452_ ;
 wire \efabless_subsystem.compute_controller_i._0455_ ;
 wire \efabless_subsystem.compute_controller_i._0457_ ;
 wire \efabless_subsystem.compute_controller_i._0458_ ;
 wire \efabless_subsystem.compute_controller_i._0460_ ;
 wire \efabless_subsystem.compute_controller_i._0461_ ;
 wire \efabless_subsystem.compute_controller_i._0462_ ;
 wire \efabless_subsystem.compute_controller_i._0463_ ;
 wire \efabless_subsystem.compute_controller_i._0464_ ;
 wire \efabless_subsystem.compute_controller_i._0465_ ;
 wire \efabless_subsystem.compute_controller_i._0466_ ;
 wire \efabless_subsystem.compute_controller_i._0467_ ;
 wire \efabless_subsystem.compute_controller_i._0468_ ;
 wire \efabless_subsystem.compute_controller_i._0469_ ;
 wire \efabless_subsystem.compute_controller_i._0470_ ;
 wire \efabless_subsystem.compute_controller_i._0471_ ;
 wire \efabless_subsystem.compute_controller_i._0472_ ;
 wire \efabless_subsystem.compute_controller_i._0473_ ;
 wire \efabless_subsystem.compute_controller_i._0474_ ;
 wire \efabless_subsystem.compute_controller_i._0475_ ;
 wire \efabless_subsystem.compute_controller_i._0476_ ;
 wire \efabless_subsystem.compute_controller_i._0477_ ;
 wire \efabless_subsystem.compute_controller_i._0478_ ;
 wire \efabless_subsystem.compute_controller_i._0479_ ;
 wire \efabless_subsystem.compute_controller_i._0480_ ;
 wire \efabless_subsystem.compute_controller_i._0481_ ;
 wire \efabless_subsystem.compute_controller_i._0482_ ;
 wire \efabless_subsystem.compute_controller_i._0483_ ;
 wire \efabless_subsystem.compute_controller_i._0484_ ;
 wire \efabless_subsystem.compute_controller_i._0485_ ;
 wire \efabless_subsystem.compute_controller_i._0486_ ;
 wire \efabless_subsystem.compute_controller_i._0487_ ;
 wire \efabless_subsystem.compute_controller_i._0488_ ;
 wire \efabless_subsystem.compute_controller_i._0489_ ;
 wire \efabless_subsystem.compute_controller_i._0490_ ;
 wire \efabless_subsystem.compute_controller_i._0491_ ;
 wire \efabless_subsystem.compute_controller_i._0492_ ;
 wire \efabless_subsystem.compute_controller_i._0493_ ;
 wire \efabless_subsystem.compute_controller_i._0494_ ;
 wire \efabless_subsystem.compute_controller_i._0495_ ;
 wire \efabless_subsystem.compute_controller_i._0496_ ;
 wire \efabless_subsystem.compute_controller_i._0497_ ;
 wire \efabless_subsystem.compute_controller_i._0498_ ;
 wire \efabless_subsystem.compute_controller_i._0499_ ;
 wire \efabless_subsystem.compute_controller_i._0500_ ;
 wire \efabless_subsystem.compute_controller_i._0501_ ;
 wire \efabless_subsystem.compute_controller_i._0502_ ;
 wire \efabless_subsystem.compute_controller_i._0503_ ;
 wire \efabless_subsystem.compute_controller_i._0504_ ;
 wire \efabless_subsystem.compute_controller_i._0505_ ;
 wire \efabless_subsystem.compute_controller_i._0506_ ;
 wire \efabless_subsystem.compute_controller_i._0507_ ;
 wire \efabless_subsystem.compute_controller_i._0508_ ;
 wire \efabless_subsystem.compute_controller_i._0509_ ;
 wire \efabless_subsystem.compute_controller_i._0510_ ;
 wire \efabless_subsystem.compute_controller_i._0511_ ;
 wire \efabless_subsystem.compute_controller_i._0512_ ;
 wire \efabless_subsystem.compute_controller_i._0513_ ;
 wire \efabless_subsystem.compute_controller_i._0514_ ;
 wire \efabless_subsystem.compute_controller_i._0515_ ;
 wire \efabless_subsystem.compute_controller_i._0516_ ;
 wire \efabless_subsystem.compute_controller_i._0517_ ;
 wire \efabless_subsystem.compute_controller_i._0518_ ;
 wire \efabless_subsystem.compute_controller_i._0519_ ;
 wire \efabless_subsystem.compute_controller_i._0520_ ;
 wire \efabless_subsystem.compute_controller_i._0521_ ;
 wire \efabless_subsystem.compute_controller_i._0522_ ;
 wire \efabless_subsystem.compute_controller_i._0523_ ;
 wire \efabless_subsystem.compute_controller_i._0524_ ;
 wire \efabless_subsystem.compute_controller_i._0525_ ;
 wire \efabless_subsystem.compute_controller_i._0526_ ;
 wire \efabless_subsystem.compute_controller_i._0527_ ;
 wire \efabless_subsystem.compute_controller_i._0528_ ;
 wire \efabless_subsystem.compute_controller_i._0529_ ;
 wire \efabless_subsystem.compute_controller_i._0530_ ;
 wire \efabless_subsystem.compute_controller_i._0531_ ;
 wire \efabless_subsystem.compute_controller_i._0532_ ;
 wire \efabless_subsystem.compute_controller_i._0533_ ;
 wire \efabless_subsystem.compute_controller_i._0534_ ;
 wire \efabless_subsystem.compute_controller_i._0535_ ;
 wire \efabless_subsystem.compute_controller_i._0536_ ;
 wire \efabless_subsystem.compute_controller_i._0537_ ;
 wire \efabless_subsystem.compute_controller_i._0538_ ;
 wire \efabless_subsystem.compute_controller_i._0539_ ;
 wire \efabless_subsystem.compute_controller_i._0540_ ;
 wire \efabless_subsystem.compute_controller_i._0541_ ;
 wire \efabless_subsystem.compute_controller_i._0542_ ;
 wire \efabless_subsystem.compute_controller_i._0543_ ;
 wire \efabless_subsystem.compute_controller_i._0544_ ;
 wire \efabless_subsystem.compute_controller_i._0545_ ;
 wire \efabless_subsystem.compute_controller_i._0546_ ;
 wire \efabless_subsystem.compute_controller_i._0547_ ;
 wire \efabless_subsystem.compute_controller_i._0548_ ;
 wire \efabless_subsystem.compute_controller_i._0549_ ;
 wire \efabless_subsystem.compute_controller_i._0550_ ;
 wire \efabless_subsystem.compute_controller_i._0551_ ;
 wire \efabless_subsystem.compute_controller_i._0552_ ;
 wire \efabless_subsystem.compute_controller_i._0553_ ;
 wire \efabless_subsystem.compute_controller_i._0554_ ;
 wire \efabless_subsystem.compute_controller_i._0555_ ;
 wire \efabless_subsystem.compute_controller_i._0556_ ;
 wire \efabless_subsystem.compute_controller_i._0557_ ;
 wire \efabless_subsystem.compute_controller_i._0558_ ;
 wire \efabless_subsystem.compute_controller_i._0559_ ;
 wire \efabless_subsystem.compute_controller_i._0560_ ;
 wire \efabless_subsystem.compute_controller_i._0561_ ;
 wire \efabless_subsystem.compute_controller_i._0562_ ;
 wire \efabless_subsystem.compute_controller_i._0563_ ;
 wire \efabless_subsystem.compute_controller_i._0564_ ;
 wire \efabless_subsystem.compute_controller_i._0565_ ;
 wire \efabless_subsystem.compute_controller_i._0566_ ;
 wire \efabless_subsystem.compute_controller_i._0567_ ;
 wire \efabless_subsystem.compute_controller_i._0568_ ;
 wire \efabless_subsystem.compute_controller_i._0569_ ;
 wire \efabless_subsystem.compute_controller_i._0570_ ;
 wire \efabless_subsystem.compute_controller_i._0571_ ;
 wire \efabless_subsystem.compute_controller_i._0572_ ;
 wire \efabless_subsystem.compute_controller_i._0573_ ;
 wire \efabless_subsystem.compute_controller_i._0574_ ;
 wire \efabless_subsystem.compute_controller_i._0575_ ;
 wire \efabless_subsystem.compute_controller_i._0576_ ;
 wire \efabless_subsystem.compute_controller_i._0577_ ;
 wire \efabless_subsystem.compute_controller_i._0578_ ;
 wire \efabless_subsystem.compute_controller_i._0579_ ;
 wire \efabless_subsystem.compute_controller_i._0580_ ;
 wire \efabless_subsystem.compute_controller_i._0581_ ;
 wire \efabless_subsystem.compute_controller_i._0582_ ;
 wire \efabless_subsystem.compute_controller_i._0583_ ;
 wire \efabless_subsystem.compute_controller_i._0584_ ;
 wire \efabless_subsystem.compute_controller_i._0585_ ;
 wire \efabless_subsystem.compute_controller_i._0586_ ;
 wire \efabless_subsystem.compute_controller_i._0587_ ;
 wire \efabless_subsystem.compute_controller_i._0588_ ;
 wire \efabless_subsystem.compute_controller_i._0589_ ;
 wire \efabless_subsystem.compute_controller_i._0590_ ;
 wire \efabless_subsystem.compute_controller_i._0591_ ;
 wire \efabless_subsystem.compute_controller_i._0592_ ;
 wire \efabless_subsystem.compute_controller_i._0593_ ;
 wire \efabless_subsystem.compute_controller_i._0594_ ;
 wire \efabless_subsystem.compute_controller_i._0595_ ;
 wire \efabless_subsystem.compute_controller_i._0596_ ;
 wire \efabless_subsystem.compute_controller_i._0597_ ;
 wire \efabless_subsystem.compute_controller_i._0598_ ;
 wire \efabless_subsystem.compute_controller_i._0599_ ;
 wire \efabless_subsystem.compute_controller_i._0600_ ;
 wire \efabless_subsystem.compute_controller_i._0601_ ;
 wire \efabless_subsystem.compute_controller_i._0602_ ;
 wire \efabless_subsystem.compute_controller_i._0603_ ;
 wire \efabless_subsystem.compute_controller_i._0604_ ;
 wire \efabless_subsystem.compute_controller_i._0605_ ;
 wire \efabless_subsystem.compute_controller_i._0606_ ;
 wire \efabless_subsystem.compute_controller_i._0607_ ;
 wire \efabless_subsystem.compute_controller_i._0608_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[0] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[10] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[11] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[12] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[13] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[14] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[15] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[1] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[2] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[3] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[4] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[5] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[6] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[7] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[8] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_d[9] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[0] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[10] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[11] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[12] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[13] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[14] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[15] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[1] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[2] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[3] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[4] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[5] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[6] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[7] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[8] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q[9] ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_edge ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg._06_ ;
 wire \efabless_subsystem.compute_controller_i.acc_done_q_reg.d ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_d ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.add_143_38.A ;
 wire \efabless_subsystem.compute_controller_i.add_143_38.Z ;
 wire \efabless_subsystem.compute_controller_i.add_157_42.Z ;
 wire \efabless_subsystem.compute_controller_i.add_163_38.A[0] ;
 wire \efabless_subsystem.compute_controller_i.add_163_38.A[1] ;
 wire \efabless_subsystem.compute_controller_i.add_163_38.Z[0] ;
 wire \efabless_subsystem.compute_controller_i.add_163_38.Z[1] ;
 wire \efabless_subsystem.compute_controller_i.add_163_38._0_ ;
 wire \efabless_subsystem.compute_controller_i.add_163_38._1_ ;
 wire \efabless_subsystem.compute_controller_i.add_163_38._2_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[0] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[10] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[11] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[12] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[13] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[14] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[15] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[1] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[2] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[3] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[4] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[5] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[6] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[7] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[8] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.A[9] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[0] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[10] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[11] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[12] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[13] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[14] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[15] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[1] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[2] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[3] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[4] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[5] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[6] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[7] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[8] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34.Z[9] ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._00_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._01_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._02_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._03_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._04_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._05_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._06_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._07_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._08_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._09_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._10_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._11_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._12_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._13_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._14_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._15_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._16_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._17_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._18_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._19_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._20_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._21_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._22_ ;
 wire \efabless_subsystem.compute_controller_i.add_175_34._23_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[0] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[10] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[11] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[12] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[13] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[14] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[15] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[1] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[2] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[3] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[4] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[5] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[6] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[7] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[8] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30.Z[9] ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._00_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._01_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._02_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._03_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._04_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._05_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._06_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._07_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._08_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._09_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._10_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._11_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._12_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._13_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._14_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._15_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._16_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._17_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._18_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._19_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._20_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._21_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._22_ ;
 wire \efabless_subsystem.compute_controller_i.add_185_30._23_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[0] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[10] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[11] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[12] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[13] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[14] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[15] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[1] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[2] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[3] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[4] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[5] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[6] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[7] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[8] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.A[9] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[0] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[10] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[11] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[12] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[13] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[14] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[15] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[1] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[2] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[3] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[4] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[5] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[6] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[7] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[8] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30.Z[9] ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._00_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._01_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._02_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._03_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._04_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._05_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._06_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._07_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._08_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._09_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._10_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._11_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._12_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._13_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._14_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._15_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._16_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._17_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._18_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._19_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._20_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._21_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._22_ ;
 wire \efabless_subsystem.compute_controller_i.add_200_30._23_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_d[1] ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_d[2] ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].d ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1].d ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8].d ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._00_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._01_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._02_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._03_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._04_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._05_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._06_ ;
 wire \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9].d ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_d[0] ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_d[1] ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].d ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1].d ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._00_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._01_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._02_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._03_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._04_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._05_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._06_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2].d ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._00_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._01_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._02_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._03_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._04_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._05_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._06_ ;
 wire \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3].d ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._07_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._08_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._09_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._10_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._11_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._12_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11._13_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[0] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[10] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[11] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[1] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[2] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[3] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[4] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[5] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[6] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[7] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[8] ;
 wire \efabless_subsystem.compute_controller_i.ctl_375_11.out_0[9] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[0] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[1] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[2] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[3] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[4] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[5] ;
 wire \efabless_subsystem.compute_controller_i.ctl_775_11.out_0[6] ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._0_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._1_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._2_ ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[0] ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[1] ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[2] ;
 wire \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[3] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[0] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[10] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[11] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[12] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[13] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[14] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[15] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[1] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[2] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[3] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[4] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[5] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[6] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[7] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[8] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_d[9] ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._06_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._00_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._01_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._02_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._03_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._04_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._05_ ;
 wire \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._06_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[0] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[10] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[11] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[12] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[13] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[14] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[15] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[1] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[2] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[3] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[4] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[5] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[6] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[7] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[8] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.A[9] ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32.Z ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._00_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._01_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._02_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._03_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._04_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._05_ ;
 wire \efabless_subsystem.compute_controller_i.gt_269_32._06_ ;
 wire \efabless_subsystem.compute_controller_i.gte_255_34.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_255_34._0_ ;
 wire \efabless_subsystem.compute_controller_i.gte_262_34.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_262_34._0_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[0] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[10] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[11] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[12] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[13] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[14] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[15] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[1] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[2] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[3] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[4] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[5] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[6] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[7] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[8] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.B[9] ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._00_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._01_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._02_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._03_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._04_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._05_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._06_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._07_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._08_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._09_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._10_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._11_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._12_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._13_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._14_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._15_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._16_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._17_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._18_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._19_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._20_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._21_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._22_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._23_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._24_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._25_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._26_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._27_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._28_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._29_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._30_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._31_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._32_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._33_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._34_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._35_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._36_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._37_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._38_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._39_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._40_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._41_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._42_ ;
 wire \efabless_subsystem.compute_controller_i.gte_286_30._43_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[0] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[10] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[11] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[12] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[13] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[14] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[15] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[16] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[17] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[18] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[19] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[1] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[20] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[21] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[22] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[23] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[24] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[25] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[26] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[27] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[28] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[29] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[2] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[30] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[31] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[3] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[4] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[5] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[6] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[7] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[8] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.B[9] ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._000_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._001_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._002_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._003_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._004_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._005_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._006_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._007_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._008_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._009_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._010_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._011_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._012_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._013_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._014_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._015_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._016_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._017_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._018_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._019_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._020_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._021_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._022_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._023_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._024_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._025_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._026_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._027_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._028_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._029_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._030_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._031_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._032_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._033_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._034_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._035_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._036_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._037_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._038_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._039_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._040_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._041_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._042_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._043_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._044_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._045_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._046_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._047_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._048_ ;
 wire \efabless_subsystem.compute_controller_i.gte_678_56._049_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[0] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[10] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[11] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[12] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[13] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[14] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[15] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[16] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[17] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[18] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[19] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[1] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[20] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[21] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[22] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[23] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[24] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[25] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[26] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[27] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[28] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[29] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[2] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[30] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[31] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[3] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[4] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[5] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[6] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[7] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[8] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.B[9] ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._000_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._001_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._002_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._003_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._004_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._005_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._006_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._007_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._008_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._009_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._010_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._011_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._012_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._013_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._014_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._015_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._016_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._017_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._018_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._019_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._020_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._021_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._022_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._023_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._024_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._025_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._026_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._027_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._028_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._029_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._030_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._031_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._032_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._033_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._034_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._035_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._036_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._037_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._038_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._039_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._040_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._041_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._042_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._043_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._044_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._045_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._046_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._047_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._048_ ;
 wire \efabless_subsystem.compute_controller_i.gte_688_48._049_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[0] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[10] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[11] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[12] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[13] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[14] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[15] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[16] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[17] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[18] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[19] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[1] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[20] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[21] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[22] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[23] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[24] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[25] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[26] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[27] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[28] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[29] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[2] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[30] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[31] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[3] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[4] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[5] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[6] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[7] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[8] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.B[9] ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._000_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._001_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._002_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._003_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._004_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._005_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._006_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._007_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._008_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._009_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._010_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._011_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._012_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._013_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._014_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._015_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._016_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._017_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._018_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._019_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._020_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._021_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._022_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._023_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._024_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._025_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._026_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._027_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._028_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._029_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._030_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._031_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._032_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._033_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._034_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._035_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._036_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._037_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._038_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._039_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._040_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._041_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._042_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._043_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._044_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._045_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._046_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._047_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._048_ ;
 wire \efabless_subsystem.compute_controller_i.gte_700_40._049_ ;
 wire \efabless_subsystem.compute_controller_i.gte_709_36.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_709_36._0_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._00_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._01_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._02_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._03_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._04_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._05_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._06_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._07_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._08_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._09_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._10_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._11_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._12_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._13_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._14_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._15_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._16_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._17_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._18_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._19_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._20_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._21_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._22_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._23_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._24_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._25_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._26_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._27_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._28_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._29_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._30_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._31_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._32_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._33_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._34_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._35_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._36_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._37_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._38_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._39_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._40_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._41_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._42_ ;
 wire \efabless_subsystem.compute_controller_i.gte_734_31._43_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31.Z ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._00_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._01_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._02_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._03_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._04_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._05_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._06_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._07_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._08_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._09_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._10_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._11_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._12_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._13_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._14_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._15_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._16_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._17_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._18_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._19_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._20_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._21_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._22_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._23_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._24_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._25_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._26_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._27_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._28_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._29_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._30_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._31_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._32_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._33_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._34_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._35_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._36_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._37_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._38_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._39_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._40_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._41_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._42_ ;
 wire \efabless_subsystem.compute_controller_i.gte_735_31._43_ ;
 wire \efabless_subsystem.compute_controller_i.i_acc_almost_done ;
 wire \efabless_subsystem.compute_controller_i.i_arr_data_valid ;
 wire \efabless_subsystem.compute_controller_i.i_start ;
 wire \efabless_subsystem.compute_controller_i.lt_156_26.Z ;
 wire \efabless_subsystem.compute_controller_i.lt_156_26._0_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35.Z ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._00_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._01_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._02_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._03_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._04_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._05_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._06_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._07_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._08_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._09_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._10_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._11_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._12_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._13_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._14_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._15_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._16_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._17_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._18_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._19_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._20_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._21_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._22_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._23_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._24_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._25_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._26_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._27_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._28_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._29_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._30_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._31_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._32_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._33_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._34_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._35_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._36_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._37_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._38_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._39_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._40_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._41_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._42_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._43_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._44_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._45_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._46_ ;
 wire \efabless_subsystem.compute_controller_i.lt_302_35._47_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g10._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g11._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g12._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g13._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g14._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g15._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g16._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g5._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g6._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g7._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g8._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g9._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_156_26.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._1_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._2_ ;
 wire \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1.z ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._1_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._2_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data3 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._1_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._2_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data3 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._1_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._2_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data3 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data4 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data5 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_749_18.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2.z ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._1_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._2_ ;
 wire \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1.z ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._08_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._09_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._10_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._11_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._12_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._13_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._14_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data4 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data5 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data7 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data8 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._08_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._09_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._10_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._11_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._12_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._13_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._14_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data4 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data5 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data7 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data8 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._08_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._09_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._10_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._11_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._12_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._13_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._14_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data4 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data5 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data7 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data8 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._00_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._01_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._02_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._03_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._04_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._05_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._06_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._07_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._08_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._09_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._10_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._11_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._12_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._13_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._14_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data3 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data4 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data5 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data7 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data8 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_269_32.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g10._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g11._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g12._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g13._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g14._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g15._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g16._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g5._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g6._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g7._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g8._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g9._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.z ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.data0 ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.data2 ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.z ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9.data1 ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9.z ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g10._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g11._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g12._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g13._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g14._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g15._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g16._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g2._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g3._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g4._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g5._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g6._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g7._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g8._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g9._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.ctl ;
 wire \efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1._0_ ;
 wire \efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1.z ;
 wire \efabless_subsystem.compute_controller_i.o_red_params_pop ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._06_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._00_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._01_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._02_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._03_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._04_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._05_ ;
 wire \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._06_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._00_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._01_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._02_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._03_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._04_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._05_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._06_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._07_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._08_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._09_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._10_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._11_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._12_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._13_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._14_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._15_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._16_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._17_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._18_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._19_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._20_ ;
 wire \efabless_subsystem.compute_controller_i.sub_302_49._21_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._00_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._01_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._02_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._03_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._04_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._05_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._06_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._07_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._08_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._09_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._10_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._11_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._12_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._13_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._14_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._15_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._16_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._17_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._18_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._19_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._20_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._21_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._22_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._23_ ;
 wire \efabless_subsystem.compute_controller_i.sub_688_68._24_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._00_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._01_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._02_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._03_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._04_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._05_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._06_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._07_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._08_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._09_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._10_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._11_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._12_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._13_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._14_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._15_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._16_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._17_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._18_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._19_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._20_ ;
 wire \efabless_subsystem.compute_controller_i.sub_700_60._21_ ;
 wire \efabless_subsystem.compute_core_i._0_ ;
 wire \efabless_subsystem.compute_core_i._1_ ;
 wire \efabless_subsystem.compute_core_i.array_acc_ready ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._000_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._002_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._003_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._137_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._138_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._139_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._140_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._141_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._142_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_ready_i ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_reg_q_reg[0][0].aclr ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._00_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._01_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._02_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._03_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._04_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._05_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._06_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0].d ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._00_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._01_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._02_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._03_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._04_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._05_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._06_ ;
 wire \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ;
 wire \efabless_subsystem.compute_core_i.fmap_reg_valid ;
 wire \efabless_subsystem.compute_core_i.i_acc_shift[0] ;
 wire \efabless_subsystem.compute_core_i.i_acc_shift[1] ;
 wire \efabless_subsystem.compute_core_i.i_acc_shift[2] ;
 wire \efabless_subsystem.compute_core_i.i_acc_shift[3] ;
 wire \efabless_subsystem.compute_core_i.i_acc_shift[4] ;
 wire \efabless_subsystem.compute_core_i.i_acc_sign ;
 wire \efabless_subsystem.compute_core_i.i_array_shftsgn[0] ;
 wire \efabless_subsystem.compute_core_i.i_array_shftsgn[1] ;
 wire \efabless_subsystem.compute_core_i.i_array_shftsgn[2] ;
 wire \efabless_subsystem.compute_core_i.i_array_shftsgn[3] ;
 wire \efabless_subsystem.compute_core_i.i_array_shftsgn_valid ;
 wire \efabless_subsystem.compute_core_i.i_fmap[0] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[10] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[11] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[12] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[13] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[14] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[15] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[16] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[17] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[18] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[19] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[1] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[20] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[21] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[22] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[23] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[24] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[25] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[26] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[27] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[28] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[29] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[2] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[30] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[31] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[32] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[33] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[34] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[35] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[36] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[37] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[38] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[39] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[3] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[40] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[41] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[42] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[43] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[44] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[45] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[46] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[47] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[48] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[49] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[4] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[50] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[51] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[52] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[53] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[54] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[55] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[56] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[57] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[58] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[59] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[5] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[60] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[61] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[62] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[63] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[6] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[7] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[8] ;
 wire \efabless_subsystem.compute_core_i.i_fmap[9] ;
 wire \efabless_subsystem.compute_core_i.i_fmap_valid ;
 wire \efabless_subsystem.compute_core_i.i_stat_cfg ;
 wire \efabless_subsystem.compute_core_i.i_weight[0] ;
 wire \efabless_subsystem.compute_core_i.i_weight[100] ;
 wire \efabless_subsystem.compute_core_i.i_weight[101] ;
 wire \efabless_subsystem.compute_core_i.i_weight[102] ;
 wire \efabless_subsystem.compute_core_i.i_weight[103] ;
 wire \efabless_subsystem.compute_core_i.i_weight[104] ;
 wire \efabless_subsystem.compute_core_i.i_weight[105] ;
 wire \efabless_subsystem.compute_core_i.i_weight[106] ;
 wire \efabless_subsystem.compute_core_i.i_weight[107] ;
 wire \efabless_subsystem.compute_core_i.i_weight[108] ;
 wire \efabless_subsystem.compute_core_i.i_weight[109] ;
 wire \efabless_subsystem.compute_core_i.i_weight[10] ;
 wire \efabless_subsystem.compute_core_i.i_weight[110] ;
 wire \efabless_subsystem.compute_core_i.i_weight[111] ;
 wire \efabless_subsystem.compute_core_i.i_weight[112] ;
 wire \efabless_subsystem.compute_core_i.i_weight[113] ;
 wire \efabless_subsystem.compute_core_i.i_weight[114] ;
 wire \efabless_subsystem.compute_core_i.i_weight[115] ;
 wire \efabless_subsystem.compute_core_i.i_weight[116] ;
 wire \efabless_subsystem.compute_core_i.i_weight[117] ;
 wire \efabless_subsystem.compute_core_i.i_weight[118] ;
 wire \efabless_subsystem.compute_core_i.i_weight[119] ;
 wire \efabless_subsystem.compute_core_i.i_weight[11] ;
 wire \efabless_subsystem.compute_core_i.i_weight[120] ;
 wire \efabless_subsystem.compute_core_i.i_weight[121] ;
 wire \efabless_subsystem.compute_core_i.i_weight[122] ;
 wire \efabless_subsystem.compute_core_i.i_weight[123] ;
 wire \efabless_subsystem.compute_core_i.i_weight[124] ;
 wire \efabless_subsystem.compute_core_i.i_weight[125] ;
 wire \efabless_subsystem.compute_core_i.i_weight[126] ;
 wire \efabless_subsystem.compute_core_i.i_weight[127] ;
 wire \efabless_subsystem.compute_core_i.i_weight[12] ;
 wire \efabless_subsystem.compute_core_i.i_weight[13] ;
 wire \efabless_subsystem.compute_core_i.i_weight[14] ;
 wire \efabless_subsystem.compute_core_i.i_weight[15] ;
 wire \efabless_subsystem.compute_core_i.i_weight[16] ;
 wire \efabless_subsystem.compute_core_i.i_weight[17] ;
 wire \efabless_subsystem.compute_core_i.i_weight[18] ;
 wire \efabless_subsystem.compute_core_i.i_weight[19] ;
 wire \efabless_subsystem.compute_core_i.i_weight[1] ;
 wire \efabless_subsystem.compute_core_i.i_weight[20] ;
 wire \efabless_subsystem.compute_core_i.i_weight[21] ;
 wire \efabless_subsystem.compute_core_i.i_weight[22] ;
 wire \efabless_subsystem.compute_core_i.i_weight[23] ;
 wire \efabless_subsystem.compute_core_i.i_weight[24] ;
 wire \efabless_subsystem.compute_core_i.i_weight[25] ;
 wire \efabless_subsystem.compute_core_i.i_weight[26] ;
 wire \efabless_subsystem.compute_core_i.i_weight[27] ;
 wire \efabless_subsystem.compute_core_i.i_weight[28] ;
 wire \efabless_subsystem.compute_core_i.i_weight[29] ;
 wire \efabless_subsystem.compute_core_i.i_weight[2] ;
 wire \efabless_subsystem.compute_core_i.i_weight[30] ;
 wire \efabless_subsystem.compute_core_i.i_weight[31] ;
 wire \efabless_subsystem.compute_core_i.i_weight[32] ;
 wire \efabless_subsystem.compute_core_i.i_weight[33] ;
 wire \efabless_subsystem.compute_core_i.i_weight[34] ;
 wire \efabless_subsystem.compute_core_i.i_weight[35] ;
 wire \efabless_subsystem.compute_core_i.i_weight[36] ;
 wire \efabless_subsystem.compute_core_i.i_weight[37] ;
 wire \efabless_subsystem.compute_core_i.i_weight[38] ;
 wire \efabless_subsystem.compute_core_i.i_weight[39] ;
 wire \efabless_subsystem.compute_core_i.i_weight[3] ;
 wire \efabless_subsystem.compute_core_i.i_weight[40] ;
 wire \efabless_subsystem.compute_core_i.i_weight[41] ;
 wire \efabless_subsystem.compute_core_i.i_weight[42] ;
 wire \efabless_subsystem.compute_core_i.i_weight[43] ;
 wire \efabless_subsystem.compute_core_i.i_weight[44] ;
 wire \efabless_subsystem.compute_core_i.i_weight[45] ;
 wire \efabless_subsystem.compute_core_i.i_weight[46] ;
 wire \efabless_subsystem.compute_core_i.i_weight[47] ;
 wire \efabless_subsystem.compute_core_i.i_weight[48] ;
 wire \efabless_subsystem.compute_core_i.i_weight[49] ;
 wire \efabless_subsystem.compute_core_i.i_weight[4] ;
 wire \efabless_subsystem.compute_core_i.i_weight[50] ;
 wire \efabless_subsystem.compute_core_i.i_weight[51] ;
 wire \efabless_subsystem.compute_core_i.i_weight[52] ;
 wire \efabless_subsystem.compute_core_i.i_weight[53] ;
 wire \efabless_subsystem.compute_core_i.i_weight[54] ;
 wire \efabless_subsystem.compute_core_i.i_weight[55] ;
 wire \efabless_subsystem.compute_core_i.i_weight[56] ;
 wire \efabless_subsystem.compute_core_i.i_weight[57] ;
 wire \efabless_subsystem.compute_core_i.i_weight[58] ;
 wire \efabless_subsystem.compute_core_i.i_weight[59] ;
 wire \efabless_subsystem.compute_core_i.i_weight[5] ;
 wire \efabless_subsystem.compute_core_i.i_weight[60] ;
 wire \efabless_subsystem.compute_core_i.i_weight[61] ;
 wire \efabless_subsystem.compute_core_i.i_weight[62] ;
 wire \efabless_subsystem.compute_core_i.i_weight[63] ;
 wire \efabless_subsystem.compute_core_i.i_weight[64] ;
 wire \efabless_subsystem.compute_core_i.i_weight[65] ;
 wire \efabless_subsystem.compute_core_i.i_weight[66] ;
 wire \efabless_subsystem.compute_core_i.i_weight[67] ;
 wire \efabless_subsystem.compute_core_i.i_weight[68] ;
 wire \efabless_subsystem.compute_core_i.i_weight[69] ;
 wire \efabless_subsystem.compute_core_i.i_weight[6] ;
 wire \efabless_subsystem.compute_core_i.i_weight[70] ;
 wire \efabless_subsystem.compute_core_i.i_weight[71] ;
 wire \efabless_subsystem.compute_core_i.i_weight[72] ;
 wire \efabless_subsystem.compute_core_i.i_weight[73] ;
 wire \efabless_subsystem.compute_core_i.i_weight[74] ;
 wire \efabless_subsystem.compute_core_i.i_weight[75] ;
 wire \efabless_subsystem.compute_core_i.i_weight[76] ;
 wire \efabless_subsystem.compute_core_i.i_weight[77] ;
 wire \efabless_subsystem.compute_core_i.i_weight[78] ;
 wire \efabless_subsystem.compute_core_i.i_weight[79] ;
 wire \efabless_subsystem.compute_core_i.i_weight[7] ;
 wire \efabless_subsystem.compute_core_i.i_weight[80] ;
 wire \efabless_subsystem.compute_core_i.i_weight[81] ;
 wire \efabless_subsystem.compute_core_i.i_weight[82] ;
 wire \efabless_subsystem.compute_core_i.i_weight[83] ;
 wire \efabless_subsystem.compute_core_i.i_weight[84] ;
 wire \efabless_subsystem.compute_core_i.i_weight[85] ;
 wire \efabless_subsystem.compute_core_i.i_weight[86] ;
 wire \efabless_subsystem.compute_core_i.i_weight[87] ;
 wire \efabless_subsystem.compute_core_i.i_weight[88] ;
 wire \efabless_subsystem.compute_core_i.i_weight[89] ;
 wire \efabless_subsystem.compute_core_i.i_weight[8] ;
 wire \efabless_subsystem.compute_core_i.i_weight[90] ;
 wire \efabless_subsystem.compute_core_i.i_weight[91] ;
 wire \efabless_subsystem.compute_core_i.i_weight[92] ;
 wire \efabless_subsystem.compute_core_i.i_weight[93] ;
 wire \efabless_subsystem.compute_core_i.i_weight[94] ;
 wire \efabless_subsystem.compute_core_i.i_weight[95] ;
 wire \efabless_subsystem.compute_core_i.i_weight[96] ;
 wire \efabless_subsystem.compute_core_i.i_weight[97] ;
 wire \efabless_subsystem.compute_core_i.i_weight[98] ;
 wire \efabless_subsystem.compute_core_i.i_weight[99] ;
 wire \efabless_subsystem.compute_core_i.i_weight[9] ;
 wire \efabless_subsystem.compute_core_i.i_weight_valid ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i._00_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i._01_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i._03_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i._04_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i._05_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i._06_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_d ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0].aclr ;
 wire \efabless_subsystem.compute_core_i.ifmap_regs_i.o_ready ;
 wire \efabless_subsystem.compute_core_i.mux_152_27.g1._0_ ;
 wire \efabless_subsystem.compute_core_i.mux_152_27.g1.data0 ;
 wire \efabless_subsystem.compute_core_i.mux_152_27.g1.data1 ;
 wire \efabless_subsystem.compute_core_i.o_array_shftsgn_ready ;
 wire \efabless_subsystem.compute_core_i.o_weight_ready ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._006_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._008_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._010_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._012_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._017_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._018_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._019_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._032_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._034_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._035_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._036_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._041_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._042_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._043_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._044_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._045_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._046_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._047_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._048_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i._049_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.acc_write_valid_reg.aclr ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.Z[0] ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.Z[1] ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._1_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._2_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._1_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._2_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_d ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1.data0 ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1.data1 ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_125_17.g1._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_132_31.g1._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1.z ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2._0_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2.z ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._00_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._01_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._02_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._03_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._04_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._05_ ;
 wire \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._06_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_reg_valid ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i._00_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i._01_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i._03_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i._04_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i._05_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i._06_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_d ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0].aclr ;
 wire \efabless_subsystem.compute_core_i.weight_reg_valid ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i._00_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i._01_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i._03_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i._04_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i._05_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i._06_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_d ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._00_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._01_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._02_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._03_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._04_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._05_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._06_ ;
 wire \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0].aclr ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED1 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED11 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED13 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED15 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED17 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED19 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED21 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED23 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED25 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED27 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED29 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED3 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED31 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED33 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED35 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED37 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED39 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED41 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED43 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED45 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED47 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED49 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED5 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED51 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED53 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED55 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED57 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED59 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED61 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED63 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED7 ;
 wire \efabless_subsystem.config_regs_i.UNCONNECTED9 ;
 wire \efabless_subsystem.config_regs_i._0000_ ;
 wire \efabless_subsystem.config_regs_i._0002_ ;
 wire \efabless_subsystem.config_regs_i._0003_ ;
 wire \efabless_subsystem.config_regs_i._0004_ ;
 wire \efabless_subsystem.config_regs_i._0005_ ;
 wire \efabless_subsystem.config_regs_i._0006_ ;
 wire \efabless_subsystem.config_regs_i._0007_ ;
 wire \efabless_subsystem.config_regs_i._0008_ ;
 wire \efabless_subsystem.config_regs_i._0009_ ;
 wire \efabless_subsystem.config_regs_i._0010_ ;
 wire \efabless_subsystem.config_regs_i._0011_ ;
 wire \efabless_subsystem.config_regs_i._0012_ ;
 wire \efabless_subsystem.config_regs_i._0013_ ;
 wire \efabless_subsystem.config_regs_i._0014_ ;
 wire \efabless_subsystem.config_regs_i._0015_ ;
 wire \efabless_subsystem.config_regs_i._0016_ ;
 wire \efabless_subsystem.config_regs_i._0017_ ;
 wire \efabless_subsystem.config_regs_i._0018_ ;
 wire \efabless_subsystem.config_regs_i._0019_ ;
 wire \efabless_subsystem.config_regs_i._0020_ ;
 wire \efabless_subsystem.config_regs_i._0021_ ;
 wire \efabless_subsystem.config_regs_i._0022_ ;
 wire \efabless_subsystem.config_regs_i._0023_ ;
 wire \efabless_subsystem.config_regs_i._0024_ ;
 wire \efabless_subsystem.config_regs_i._0025_ ;
 wire \efabless_subsystem.config_regs_i._0026_ ;
 wire \efabless_subsystem.config_regs_i._0027_ ;
 wire \efabless_subsystem.config_regs_i._0028_ ;
 wire \efabless_subsystem.config_regs_i._0029_ ;
 wire \efabless_subsystem.config_regs_i._0030_ ;
 wire \efabless_subsystem.config_regs_i._0031_ ;
 wire \efabless_subsystem.config_regs_i._0032_ ;
 wire \efabless_subsystem.config_regs_i._0033_ ;
 wire \efabless_subsystem.config_regs_i._0034_ ;
 wire \efabless_subsystem.config_regs_i._0035_ ;
 wire \efabless_subsystem.config_regs_i._0036_ ;
 wire \efabless_subsystem.config_regs_i._0037_ ;
 wire \efabless_subsystem.config_regs_i._0038_ ;
 wire \efabless_subsystem.config_regs_i._0039_ ;
 wire \efabless_subsystem.config_regs_i._0040_ ;
 wire \efabless_subsystem.config_regs_i._0041_ ;
 wire \efabless_subsystem.config_regs_i._0044_ ;
 wire \efabless_subsystem.config_regs_i._0078_ ;
 wire \efabless_subsystem.config_regs_i._0079_ ;
 wire \efabless_subsystem.config_regs_i._0080_ ;
 wire \efabless_subsystem.config_regs_i._0083_ ;
 wire \efabless_subsystem.config_regs_i._0084_ ;
 wire \efabless_subsystem.config_regs_i._0085_ ;
 wire \efabless_subsystem.config_regs_i._0086_ ;
 wire \efabless_subsystem.config_regs_i._0090_ ;
 wire \efabless_subsystem.config_regs_i._0092_ ;
 wire \efabless_subsystem.config_regs_i._0093_ ;
 wire \efabless_subsystem.config_regs_i._0094_ ;
 wire \efabless_subsystem.config_regs_i._0095_ ;
 wire \efabless_subsystem.config_regs_i._0096_ ;
 wire \efabless_subsystem.config_regs_i._0097_ ;
 wire \efabless_subsystem.config_regs_i._0098_ ;
 wire \efabless_subsystem.config_regs_i._0099_ ;
 wire \efabless_subsystem.config_regs_i._0100_ ;
 wire \efabless_subsystem.config_regs_i._0101_ ;
 wire \efabless_subsystem.config_regs_i._0102_ ;
 wire \efabless_subsystem.config_regs_i._0103_ ;
 wire \efabless_subsystem.config_regs_i._0104_ ;
 wire \efabless_subsystem.config_regs_i._0105_ ;
 wire \efabless_subsystem.config_regs_i._0106_ ;
 wire \efabless_subsystem.config_regs_i._0107_ ;
 wire \efabless_subsystem.config_regs_i._0108_ ;
 wire \efabless_subsystem.config_regs_i._0109_ ;
 wire \efabless_subsystem.config_regs_i._0110_ ;
 wire \efabless_subsystem.config_regs_i._0111_ ;
 wire \efabless_subsystem.config_regs_i._0112_ ;
 wire \efabless_subsystem.config_regs_i._0113_ ;
 wire \efabless_subsystem.config_regs_i._0114_ ;
 wire \efabless_subsystem.config_regs_i._0115_ ;
 wire \efabless_subsystem.config_regs_i._0116_ ;
 wire \efabless_subsystem.config_regs_i._0117_ ;
 wire \efabless_subsystem.config_regs_i._0118_ ;
 wire \efabless_subsystem.config_regs_i._0119_ ;
 wire \efabless_subsystem.config_regs_i._0120_ ;
 wire \efabless_subsystem.config_regs_i._0121_ ;
 wire \efabless_subsystem.config_regs_i._0122_ ;
 wire \efabless_subsystem.config_regs_i._0123_ ;
 wire \efabless_subsystem.config_regs_i._0124_ ;
 wire \efabless_subsystem.config_regs_i._0125_ ;
 wire \efabless_subsystem.config_regs_i._0126_ ;
 wire \efabless_subsystem.config_regs_i._0127_ ;
 wire \efabless_subsystem.config_regs_i._0159_ ;
 wire \efabless_subsystem.config_regs_i._0160_ ;
 wire \efabless_subsystem.config_regs_i._0161_ ;
 wire \efabless_subsystem.config_regs_i._0162_ ;
 wire \efabless_subsystem.config_regs_i._0170_ ;
 wire \efabless_subsystem.config_regs_i._0181_ ;
 wire \efabless_subsystem.config_regs_i._0184_ ;
 wire \efabless_subsystem.config_regs_i._0185_ ;
 wire \efabless_subsystem.config_regs_i._0186_ ;
 wire \efabless_subsystem.config_regs_i._0187_ ;
 wire \efabless_subsystem.config_regs_i._0188_ ;
 wire \efabless_subsystem.config_regs_i._0189_ ;
 wire \efabless_subsystem.config_regs_i._0190_ ;
 wire \efabless_subsystem.config_regs_i._0191_ ;
 wire \efabless_subsystem.config_regs_i._0192_ ;
 wire \efabless_subsystem.config_regs_i._0193_ ;
 wire \efabless_subsystem.config_regs_i._0194_ ;
 wire \efabless_subsystem.config_regs_i._0202_ ;
 wire \efabless_subsystem.config_regs_i._0213_ ;
 wire \efabless_subsystem.config_regs_i._0216_ ;
 wire \efabless_subsystem.config_regs_i._0217_ ;
 wire \efabless_subsystem.config_regs_i._0218_ ;
 wire \efabless_subsystem.config_regs_i._0219_ ;
 wire \efabless_subsystem.config_regs_i._0220_ ;
 wire \efabless_subsystem.config_regs_i._0221_ ;
 wire \efabless_subsystem.config_regs_i._0222_ ;
 wire \efabless_subsystem.config_regs_i._0223_ ;
 wire \efabless_subsystem.config_regs_i._0234_ ;
 wire \efabless_subsystem.config_regs_i._0245_ ;
 wire \efabless_subsystem.config_regs_i._0248_ ;
 wire \efabless_subsystem.config_regs_i._0249_ ;
 wire \efabless_subsystem.config_regs_i._0250_ ;
 wire \efabless_subsystem.config_regs_i._0251_ ;
 wire \efabless_subsystem.config_regs_i._0252_ ;
 wire \efabless_subsystem.config_regs_i._0253_ ;
 wire \efabless_subsystem.config_regs_i._0255_ ;
 wire \efabless_subsystem.config_regs_i._0266_ ;
 wire \efabless_subsystem.config_regs_i._0277_ ;
 wire \efabless_subsystem.config_regs_i._0280_ ;
 wire \efabless_subsystem.config_regs_i._0281_ ;
 wire \efabless_subsystem.config_regs_i._0282_ ;
 wire \efabless_subsystem.config_regs_i._0283_ ;
 wire \efabless_subsystem.config_regs_i._0284_ ;
 wire \efabless_subsystem.config_regs_i._0285_ ;
 wire \efabless_subsystem.config_regs_i._0351_ ;
 wire \efabless_subsystem.config_regs_i._0352_ ;
 wire \efabless_subsystem.config_regs_i._0385_ ;
 wire \efabless_subsystem.config_regs_i._0386_ ;
 wire \efabless_subsystem.config_regs_i._0419_ ;
 wire \efabless_subsystem.config_regs_i._0420_ ;
 wire \efabless_subsystem.config_regs_i._0421_ ;
 wire \efabless_subsystem.config_regs_i._0519_ ;
 wire \efabless_subsystem.config_regs_i._0520_ ;
 wire \efabless_subsystem.config_regs_i._0521_ ;
 wire \efabless_subsystem.config_regs_i._0522_ ;
 wire \efabless_subsystem.config_regs_i._0524_ ;
 wire \efabless_subsystem.config_regs_i._0525_ ;
 wire \efabless_subsystem.config_regs_i._0526_ ;
 wire \efabless_subsystem.config_regs_i._0527_ ;
 wire \efabless_subsystem.config_regs_i._0528_ ;
 wire \efabless_subsystem.config_regs_i._0529_ ;
 wire \efabless_subsystem.config_regs_i._0530_ ;
 wire \efabless_subsystem.config_regs_i._0531_ ;
 wire \efabless_subsystem.config_regs_i._0532_ ;
 wire \efabless_subsystem.config_regs_i._0533_ ;
 wire \efabless_subsystem.config_regs_i._0536_ ;
 wire \efabless_subsystem.config_regs_i._0569_ ;
 wire \efabless_subsystem.config_regs_i._0570_ ;
 wire \efabless_subsystem.config_regs_i._0571_ ;
 wire \efabless_subsystem.config_regs_i._0572_ ;
 wire \efabless_subsystem.config_regs_i._0819_ ;
 wire \efabless_subsystem.config_regs_i._0820_ ;
 wire \efabless_subsystem.config_regs_i._0821_ ;
 wire \efabless_subsystem.config_regs_i._0854_ ;
 wire \efabless_subsystem.config_regs_i._0855_ ;
 wire \efabless_subsystem.config_regs_i._0856_ ;
 wire \efabless_subsystem.config_regs_i._0953_ ;
 wire \efabless_subsystem.config_regs_i._0954_ ;
 wire \efabless_subsystem.config_regs_i._0955_ ;
 wire \efabless_subsystem.config_regs_i._0956_ ;
 wire \efabless_subsystem.config_regs_i._0957_ ;
 wire \efabless_subsystem.config_regs_i._0958_ ;
 wire \efabless_subsystem.config_regs_i._0959_ ;
 wire \efabless_subsystem.config_regs_i._0960_ ;
 wire \efabless_subsystem.config_regs_i._0961_ ;
 wire \efabless_subsystem.config_regs_i._0962_ ;
 wire \efabless_subsystem.config_regs_i._0963_ ;
 wire \efabless_subsystem.config_regs_i._0964_ ;
 wire \efabless_subsystem.config_regs_i._0965_ ;
 wire \efabless_subsystem.config_regs_i._0966_ ;
 wire \efabless_subsystem.config_regs_i._0967_ ;
 wire \efabless_subsystem.config_regs_i._0968_ ;
 wire \efabless_subsystem.config_regs_i._0969_ ;
 wire \efabless_subsystem.config_regs_i._0970_ ;
 wire \efabless_subsystem.config_regs_i._0971_ ;
 wire \efabless_subsystem.config_regs_i._0972_ ;
 wire \efabless_subsystem.config_regs_i._0973_ ;
 wire \efabless_subsystem.config_regs_i._0974_ ;
 wire \efabless_subsystem.config_regs_i._0975_ ;
 wire \efabless_subsystem.config_regs_i._0976_ ;
 wire \efabless_subsystem.config_regs_i._0977_ ;
 wire \efabless_subsystem.config_regs_i._0978_ ;
 wire \efabless_subsystem.config_regs_i._0979_ ;
 wire \efabless_subsystem.config_regs_i._0980_ ;
 wire \efabless_subsystem.config_regs_i._0981_ ;
 wire \efabless_subsystem.config_regs_i._0982_ ;
 wire \efabless_subsystem.config_regs_i._0983_ ;
 wire \efabless_subsystem.config_regs_i._0984_ ;
 wire \efabless_subsystem.config_regs_i._0985_ ;
 wire \efabless_subsystem.config_regs_i._0986_ ;
 wire \efabless_subsystem.config_regs_i._0987_ ;
 wire \efabless_subsystem.config_regs_i._0988_ ;
 wire \efabless_subsystem.config_regs_i._0989_ ;
 wire \efabless_subsystem.config_regs_i._0990_ ;
 wire \efabless_subsystem.config_regs_i._0991_ ;
 wire \efabless_subsystem.config_regs_i._0992_ ;
 wire \efabless_subsystem.config_regs_i._0993_ ;
 wire \efabless_subsystem.config_regs_i._0994_ ;
 wire \efabless_subsystem.config_regs_i._0995_ ;
 wire \efabless_subsystem.config_regs_i._0996_ ;
 wire \efabless_subsystem.config_regs_i._0997_ ;
 wire \efabless_subsystem.config_regs_i._0998_ ;
 wire \efabless_subsystem.config_regs_i._0999_ ;
 wire \efabless_subsystem.config_regs_i._1000_ ;
 wire \efabless_subsystem.config_regs_i._1001_ ;
 wire \efabless_subsystem.config_regs_i._1002_ ;
 wire \efabless_subsystem.config_regs_i._1003_ ;
 wire \efabless_subsystem.config_regs_i._1004_ ;
 wire \efabless_subsystem.config_regs_i._1005_ ;
 wire \efabless_subsystem.config_regs_i._1006_ ;
 wire \efabless_subsystem.config_regs_i._1007_ ;
 wire \efabless_subsystem.config_regs_i._1008_ ;
 wire \efabless_subsystem.config_regs_i._1009_ ;
 wire \efabless_subsystem.config_regs_i._1010_ ;
 wire \efabless_subsystem.config_regs_i._1011_ ;
 wire \efabless_subsystem.config_regs_i._1012_ ;
 wire \efabless_subsystem.config_regs_i._1013_ ;
 wire \efabless_subsystem.config_regs_i._1014_ ;
 wire \efabless_subsystem.config_regs_i._1015_ ;
 wire \efabless_subsystem.config_regs_i._1016_ ;
 wire \efabless_subsystem.config_regs_i._1017_ ;
 wire \efabless_subsystem.config_regs_i._1018_ ;
 wire \efabless_subsystem.config_regs_i._1019_ ;
 wire \efabless_subsystem.config_regs_i._1020_ ;
 wire \efabless_subsystem.config_regs_i._1021_ ;
 wire \efabless_subsystem.config_regs_i._1022_ ;
 wire \efabless_subsystem.config_regs_i._1023_ ;
 wire \efabless_subsystem.config_regs_i._1024_ ;
 wire \efabless_subsystem.config_regs_i._1025_ ;
 wire \efabless_subsystem.config_regs_i._1026_ ;
 wire \efabless_subsystem.config_regs_i._1027_ ;
 wire \efabless_subsystem.config_regs_i._1028_ ;
 wire \efabless_subsystem.config_regs_i._1029_ ;
 wire \efabless_subsystem.config_regs_i._1030_ ;
 wire \efabless_subsystem.config_regs_i._1031_ ;
 wire \efabless_subsystem.config_regs_i._1032_ ;
 wire \efabless_subsystem.config_regs_i._1033_ ;
 wire \efabless_subsystem.config_regs_i._1034_ ;
 wire \efabless_subsystem.config_regs_i._1035_ ;
 wire \efabless_subsystem.config_regs_i._1036_ ;
 wire \efabless_subsystem.config_regs_i._1037_ ;
 wire \efabless_subsystem.config_regs_i._1038_ ;
 wire \efabless_subsystem.config_regs_i._1039_ ;
 wire \efabless_subsystem.config_regs_i._1040_ ;
 wire \efabless_subsystem.config_regs_i._1041_ ;
 wire \efabless_subsystem.config_regs_i._1042_ ;
 wire \efabless_subsystem.config_regs_i._1043_ ;
 wire \efabless_subsystem.config_regs_i._1044_ ;
 wire \efabless_subsystem.config_regs_i._1045_ ;
 wire \efabless_subsystem.config_regs_i._1046_ ;
 wire \efabless_subsystem.config_regs_i._1047_ ;
 wire \efabless_subsystem.config_regs_i._1048_ ;
 wire \efabless_subsystem.config_regs_i._1049_ ;
 wire \efabless_subsystem.config_regs_i._1050_ ;
 wire \efabless_subsystem.config_regs_i._1051_ ;
 wire \efabless_subsystem.config_regs_i._1052_ ;
 wire \efabless_subsystem.config_regs_i._1053_ ;
 wire \efabless_subsystem.config_regs_i._1054_ ;
 wire \efabless_subsystem.config_regs_i._1055_ ;
 wire \efabless_subsystem.config_regs_i._1056_ ;
 wire \efabless_subsystem.config_regs_i._1057_ ;
 wire \efabless_subsystem.config_regs_i._1058_ ;
 wire \efabless_subsystem.config_regs_i._1059_ ;
 wire \efabless_subsystem.config_regs_i._1060_ ;
 wire \efabless_subsystem.config_regs_i._1061_ ;
 wire \efabless_subsystem.config_regs_i._1062_ ;
 wire \efabless_subsystem.config_regs_i._1063_ ;
 wire \efabless_subsystem.config_regs_i._1064_ ;
 wire \efabless_subsystem.config_regs_i._1065_ ;
 wire \efabless_subsystem.config_regs_i._1066_ ;
 wire \efabless_subsystem.config_regs_i._1067_ ;
 wire \efabless_subsystem.config_regs_i._1068_ ;
 wire \efabless_subsystem.config_regs_i._1069_ ;
 wire \efabless_subsystem.config_regs_i._1070_ ;
 wire \efabless_subsystem.config_regs_i._1071_ ;
 wire \efabless_subsystem.config_regs_i._1072_ ;
 wire \efabless_subsystem.config_regs_i._1073_ ;
 wire \efabless_subsystem.config_regs_i._1074_ ;
 wire \efabless_subsystem.config_regs_i._1075_ ;
 wire \efabless_subsystem.config_regs_i._1076_ ;
 wire \efabless_subsystem.config_regs_i._1077_ ;
 wire \efabless_subsystem.config_regs_i._1078_ ;
 wire \efabless_subsystem.config_regs_i._1079_ ;
 wire \efabless_subsystem.config_regs_i._1080_ ;
 wire \efabless_subsystem.config_regs_i._1081_ ;
 wire \efabless_subsystem.config_regs_i._1082_ ;
 wire \efabless_subsystem.config_regs_i._1083_ ;
 wire \efabless_subsystem.config_regs_i._1084_ ;
 wire \efabless_subsystem.config_regs_i._1085_ ;
 wire \efabless_subsystem.config_regs_i._1086_ ;
 wire \efabless_subsystem.config_regs_i._1087_ ;
 wire \efabless_subsystem.config_regs_i._1088_ ;
 wire \efabless_subsystem.config_regs_i._1089_ ;
 wire \efabless_subsystem.config_regs_i._1090_ ;
 wire \efabless_subsystem.config_regs_i._1091_ ;
 wire \efabless_subsystem.config_regs_i._1092_ ;
 wire \efabless_subsystem.config_regs_i._1093_ ;
 wire \efabless_subsystem.config_regs_i._1094_ ;
 wire \efabless_subsystem.config_regs_i._1095_ ;
 wire \efabless_subsystem.config_regs_i._1096_ ;
 wire \efabless_subsystem.config_regs_i._1097_ ;
 wire \efabless_subsystem.config_regs_i._1098_ ;
 wire \efabless_subsystem.config_regs_i._1099_ ;
 wire \efabless_subsystem.config_regs_i._1100_ ;
 wire \efabless_subsystem.config_regs_i._1101_ ;
 wire \efabless_subsystem.config_regs_i._1102_ ;
 wire \efabless_subsystem.config_regs_i._1103_ ;
 wire \efabless_subsystem.config_regs_i._1104_ ;
 wire \efabless_subsystem.config_regs_i._1105_ ;
 wire \efabless_subsystem.config_regs_i._1106_ ;
 wire \efabless_subsystem.config_regs_i._1107_ ;
 wire \efabless_subsystem.config_regs_i._1108_ ;
 wire \efabless_subsystem.config_regs_i._1109_ ;
 wire \efabless_subsystem.config_regs_i._1110_ ;
 wire \efabless_subsystem.config_regs_i._1111_ ;
 wire \efabless_subsystem.config_regs_i._1112_ ;
 wire \efabless_subsystem.config_regs_i._1113_ ;
 wire \efabless_subsystem.config_regs_i._1114_ ;
 wire \efabless_subsystem.config_regs_i._1115_ ;
 wire \efabless_subsystem.config_regs_i._1116_ ;
 wire \efabless_subsystem.config_regs_i._1117_ ;
 wire \efabless_subsystem.config_regs_i._1118_ ;
 wire \efabless_subsystem.config_regs_i._1119_ ;
 wire \efabless_subsystem.config_regs_i._1120_ ;
 wire \efabless_subsystem.config_regs_i._1121_ ;
 wire \efabless_subsystem.config_regs_i._1122_ ;
 wire \efabless_subsystem.config_regs_i._1123_ ;
 wire \efabless_subsystem.config_regs_i._1124_ ;
 wire \efabless_subsystem.config_regs_i._1125_ ;
 wire \efabless_subsystem.config_regs_i._1126_ ;
 wire \efabless_subsystem.config_regs_i._1127_ ;
 wire \efabless_subsystem.config_regs_i._1128_ ;
 wire \efabless_subsystem.config_regs_i._1129_ ;
 wire \efabless_subsystem.config_regs_i._1130_ ;
 wire \efabless_subsystem.config_regs_i._1131_ ;
 wire \efabless_subsystem.config_regs_i._1132_ ;
 wire \efabless_subsystem.config_regs_i._1133_ ;
 wire \efabless_subsystem.config_regs_i._1134_ ;
 wire \efabless_subsystem.config_regs_i._1135_ ;
 wire \efabless_subsystem.config_regs_i._1136_ ;
 wire \efabless_subsystem.config_regs_i._1137_ ;
 wire \efabless_subsystem.config_regs_i._1138_ ;
 wire \efabless_subsystem.config_regs_i._1139_ ;
 wire \efabless_subsystem.config_regs_i._1140_ ;
 wire \efabless_subsystem.config_regs_i._1141_ ;
 wire \efabless_subsystem.config_regs_i._1142_ ;
 wire \efabless_subsystem.config_regs_i._1143_ ;
 wire \efabless_subsystem.config_regs_i._1144_ ;
 wire \efabless_subsystem.config_regs_i._1145_ ;
 wire \efabless_subsystem.config_regs_i._1146_ ;
 wire \efabless_subsystem.config_regs_i._1147_ ;
 wire \efabless_subsystem.config_regs_i._1148_ ;
 wire \efabless_subsystem.config_regs_i._1149_ ;
 wire \efabless_subsystem.config_regs_i._1150_ ;
 wire \efabless_subsystem.config_regs_i._1151_ ;
 wire \efabless_subsystem.config_regs_i._1245_ ;
 wire \efabless_subsystem.config_regs_i._1246_ ;
 wire \efabless_subsystem.config_regs_i._1247_ ;
 wire \efabless_subsystem.config_regs_i._1248_ ;
 wire \efabless_subsystem.config_regs_i._1249_ ;
 wire \efabless_subsystem.config_regs_i._1250_ ;
 wire \efabless_subsystem.config_regs_i._1251_ ;
 wire \efabless_subsystem.config_regs_i._1252_ ;
 wire \efabless_subsystem.config_regs_i._1253_ ;
 wire \efabless_subsystem.config_regs_i._1254_ ;
 wire \efabless_subsystem.config_regs_i._1255_ ;
 wire \efabless_subsystem.config_regs_i._1256_ ;
 wire \efabless_subsystem.config_regs_i._1278_ ;
 wire \efabless_subsystem.config_regs_i._1279_ ;
 wire \efabless_subsystem.config_regs_i._1280_ ;
 wire \efabless_subsystem.config_regs_i._1311_ ;
 wire \efabless_subsystem.config_regs_i._1312_ ;
 wire \efabless_subsystem.config_regs_i._1313_ ;
 wire \efabless_subsystem.config_regs_i._1320_ ;
 wire \efabless_subsystem.config_regs_i._1321_ ;
 wire \efabless_subsystem.config_regs_i._1322_ ;
 wire \efabless_subsystem.config_regs_i._1323_ ;
 wire \efabless_subsystem.config_regs_i._1324_ ;
 wire \efabless_subsystem.config_regs_i._1325_ ;
 wire \efabless_subsystem.config_regs_i._1326_ ;
 wire \efabless_subsystem.config_regs_i._1327_ ;
 wire \efabless_subsystem.config_regs_i._1328_ ;
 wire \efabless_subsystem.config_regs_i._1329_ ;
 wire \efabless_subsystem.config_regs_i._1330_ ;
 wire \efabless_subsystem.config_regs_i._1331_ ;
 wire \efabless_subsystem.config_regs_i._1332_ ;
 wire \efabless_subsystem.config_regs_i._1333_ ;
 wire \efabless_subsystem.config_regs_i._1334_ ;
 wire \efabless_subsystem.config_regs_i._1335_ ;
 wire \efabless_subsystem.config_regs_i._1336_ ;
 wire \efabless_subsystem.config_regs_i._1337_ ;
 wire \efabless_subsystem.config_regs_i._1338_ ;
 wire \efabless_subsystem.config_regs_i._1339_ ;
 wire \efabless_subsystem.config_regs_i._1340_ ;
 wire \efabless_subsystem.config_regs_i._1341_ ;
 wire \efabless_subsystem.config_regs_i._1342_ ;
 wire \efabless_subsystem.config_regs_i._1343_ ;
 wire \efabless_subsystem.config_regs_i._1344_ ;
 wire \efabless_subsystem.config_regs_i._1345_ ;
 wire \efabless_subsystem.config_regs_i._1346_ ;
 wire \efabless_subsystem.config_regs_i._1347_ ;
 wire \efabless_subsystem.config_regs_i._1348_ ;
 wire \efabless_subsystem.config_regs_i._1349_ ;
 wire \efabless_subsystem.config_regs_i._1350_ ;
 wire \efabless_subsystem.config_regs_i._1351_ ;
 wire \efabless_subsystem.config_regs_i._1352_ ;
 wire \efabless_subsystem.config_regs_i._1374_ ;
 wire \efabless_subsystem.config_regs_i._1375_ ;
 wire \efabless_subsystem.config_regs_i._1376_ ;
 wire \efabless_subsystem.config_regs_i._1407_ ;
 wire \efabless_subsystem.config_regs_i._1408_ ;
 wire \efabless_subsystem.config_regs_i._1409_ ;
 wire \efabless_subsystem.config_regs_i._1416_ ;
 wire \efabless_subsystem.config_regs_i._1417_ ;
 wire \efabless_subsystem.config_regs_i._1418_ ;
 wire \efabless_subsystem.config_regs_i._1419_ ;
 wire \efabless_subsystem.config_regs_i._1420_ ;
 wire \efabless_subsystem.config_regs_i._1421_ ;
 wire \efabless_subsystem.config_regs_i._1422_ ;
 wire \efabless_subsystem.config_regs_i._1423_ ;
 wire \efabless_subsystem.config_regs_i._1424_ ;
 wire \efabless_subsystem.config_regs_i._1425_ ;
 wire \efabless_subsystem.config_regs_i._1426_ ;
 wire \efabless_subsystem.config_regs_i._1427_ ;
 wire \efabless_subsystem.config_regs_i._1428_ ;
 wire \efabless_subsystem.config_regs_i._1429_ ;
 wire \efabless_subsystem.config_regs_i._1430_ ;
 wire \efabless_subsystem.config_regs_i._1431_ ;
 wire \efabless_subsystem.config_regs_i._1432_ ;
 wire \efabless_subsystem.config_regs_i._1433_ ;
 wire \efabless_subsystem.config_regs_i._1434_ ;
 wire \efabless_subsystem.config_regs_i._1435_ ;
 wire \efabless_subsystem.config_regs_i._1436_ ;
 wire \efabless_subsystem.config_regs_i._1437_ ;
 wire \efabless_subsystem.config_regs_i._1438_ ;
 wire \efabless_subsystem.config_regs_i._1439_ ;
 wire \efabless_subsystem.config_regs_i._1470_ ;
 wire \efabless_subsystem.config_regs_i._1471_ ;
 wire \efabless_subsystem.config_regs_i._1472_ ;
 wire \efabless_subsystem.config_regs_i._1503_ ;
 wire \efabless_subsystem.config_regs_i._1504_ ;
 wire \efabless_subsystem.config_regs_i._1505_ ;
 wire \efabless_subsystem.config_regs_i._1512_ ;
 wire \efabless_subsystem.config_regs_i._1513_ ;
 wire \efabless_subsystem.config_regs_i._1514_ ;
 wire \efabless_subsystem.config_regs_i._1515_ ;
 wire \efabless_subsystem.config_regs_i._1516_ ;
 wire \efabless_subsystem.config_regs_i._1517_ ;
 wire \efabless_subsystem.config_regs_i._1518_ ;
 wire \efabless_subsystem.config_regs_i._1519_ ;
 wire \efabless_subsystem.config_regs_i._1520_ ;
 wire \efabless_subsystem.config_regs_i._1521_ ;
 wire \efabless_subsystem.config_regs_i._1522_ ;
 wire \efabless_subsystem.config_regs_i._1523_ ;
 wire \efabless_subsystem.config_regs_i._1524_ ;
 wire \efabless_subsystem.config_regs_i._1525_ ;
 wire \efabless_subsystem.config_regs_i._1526_ ;
 wire \efabless_subsystem.config_regs_i._1527_ ;
 wire \efabless_subsystem.config_regs_i._1528_ ;
 wire \efabless_subsystem.config_regs_i._1529_ ;
 wire \efabless_subsystem.config_regs_i._1533_ ;
 wire \efabless_subsystem.config_regs_i._1534_ ;
 wire \efabless_subsystem.config_regs_i._1535_ ;
 wire \efabless_subsystem.config_regs_i._1566_ ;
 wire \efabless_subsystem.config_regs_i._1567_ ;
 wire \efabless_subsystem.config_regs_i._1568_ ;
 wire \efabless_subsystem.config_regs_i._1599_ ;
 wire \efabless_subsystem.config_regs_i._1600_ ;
 wire \efabless_subsystem.config_regs_i._1601_ ;
 wire \efabless_subsystem.config_regs_i._1608_ ;
 wire \efabless_subsystem.config_regs_i._1609_ ;
 wire \efabless_subsystem.config_regs_i._1610_ ;
 wire \efabless_subsystem.config_regs_i._1611_ ;
 wire \efabless_subsystem.config_regs_i._1612_ ;
 wire \efabless_subsystem.config_regs_i._1613_ ;
 wire \efabless_subsystem.config_regs_i._1614_ ;
 wire \efabless_subsystem.config_regs_i._1615_ ;
 wire \efabless_subsystem.config_regs_i._1616_ ;
 wire \efabless_subsystem.config_regs_i._1617_ ;
 wire \efabless_subsystem.config_regs_i._1618_ ;
 wire \efabless_subsystem.config_regs_i._1619_ ;
 wire \efabless_subsystem.config_regs_i._1620_ ;
 wire \efabless_subsystem.config_regs_i._1621_ ;
 wire \efabless_subsystem.config_regs_i._1622_ ;
 wire \efabless_subsystem.config_regs_i._1623_ ;
 wire \efabless_subsystem.config_regs_i._1624_ ;
 wire \efabless_subsystem.config_regs_i._1625_ ;
 wire \efabless_subsystem.config_regs_i._1821_ ;
 wire \efabless_subsystem.config_regs_i._1822_ ;
 wire \efabless_subsystem.config_regs_i._1823_ ;
 wire \efabless_subsystem.config_regs_i._1824_ ;
 wire \efabless_subsystem.config_regs_i._1825_ ;
 wire \efabless_subsystem.config_regs_i._1826_ ;
 wire \efabless_subsystem.config_regs_i._1827_ ;
 wire \efabless_subsystem.config_regs_i._1828_ ;
 wire \efabless_subsystem.config_regs_i._1829_ ;
 wire \efabless_subsystem.config_regs_i._1830_ ;
 wire \efabless_subsystem.config_regs_i._1831_ ;
 wire \efabless_subsystem.config_regs_i._1832_ ;
 wire \efabless_subsystem.config_regs_i._1854_ ;
 wire \efabless_subsystem.config_regs_i._1855_ ;
 wire \efabless_subsystem.config_regs_i._1856_ ;
 wire \efabless_subsystem.config_regs_i._1887_ ;
 wire \efabless_subsystem.config_regs_i._1888_ ;
 wire \efabless_subsystem.config_regs_i._1889_ ;
 wire \efabless_subsystem.config_regs_i._1896_ ;
 wire \efabless_subsystem.config_regs_i._1897_ ;
 wire \efabless_subsystem.config_regs_i._1898_ ;
 wire \efabless_subsystem.config_regs_i._1899_ ;
 wire \efabless_subsystem.config_regs_i._1900_ ;
 wire \efabless_subsystem.config_regs_i._1901_ ;
 wire \efabless_subsystem.config_regs_i._1902_ ;
 wire \efabless_subsystem.config_regs_i._1903_ ;
 wire \efabless_subsystem.config_regs_i._1904_ ;
 wire \efabless_subsystem.config_regs_i._1905_ ;
 wire \efabless_subsystem.config_regs_i._1906_ ;
 wire \efabless_subsystem.config_regs_i._1907_ ;
 wire \efabless_subsystem.config_regs_i._1908_ ;
 wire \efabless_subsystem.config_regs_i._1909_ ;
 wire \efabless_subsystem.config_regs_i._1910_ ;
 wire \efabless_subsystem.config_regs_i._1911_ ;
 wire \efabless_subsystem.config_regs_i._1912_ ;
 wire \efabless_subsystem.config_regs_i._1913_ ;
 wire \efabless_subsystem.config_regs_i._1914_ ;
 wire \efabless_subsystem.config_regs_i._1915_ ;
 wire \efabless_subsystem.config_regs_i._1916_ ;
 wire \efabless_subsystem.config_regs_i._1917_ ;
 wire \efabless_subsystem.config_regs_i._1918_ ;
 wire \efabless_subsystem.config_regs_i._1919_ ;
 wire \efabless_subsystem.config_regs_i._1920_ ;
 wire \efabless_subsystem.config_regs_i._1921_ ;
 wire \efabless_subsystem.config_regs_i._1922_ ;
 wire \efabless_subsystem.config_regs_i._1923_ ;
 wire \efabless_subsystem.config_regs_i._1924_ ;
 wire \efabless_subsystem.config_regs_i._1925_ ;
 wire \efabless_subsystem.config_regs_i._1926_ ;
 wire \efabless_subsystem.config_regs_i._1927_ ;
 wire \efabless_subsystem.config_regs_i._1928_ ;
 wire \efabless_subsystem.config_regs_i._1950_ ;
 wire \efabless_subsystem.config_regs_i._1951_ ;
 wire \efabless_subsystem.config_regs_i._1952_ ;
 wire \efabless_subsystem.config_regs_i._1983_ ;
 wire \efabless_subsystem.config_regs_i._1984_ ;
 wire \efabless_subsystem.config_regs_i._1985_ ;
 wire \efabless_subsystem.config_regs_i._1992_ ;
 wire \efabless_subsystem.config_regs_i._1993_ ;
 wire \efabless_subsystem.config_regs_i._1994_ ;
 wire \efabless_subsystem.config_regs_i._1995_ ;
 wire \efabless_subsystem.config_regs_i._1996_ ;
 wire \efabless_subsystem.config_regs_i._1997_ ;
 wire \efabless_subsystem.config_regs_i._1998_ ;
 wire \efabless_subsystem.config_regs_i._1999_ ;
 wire \efabless_subsystem.config_regs_i._2000_ ;
 wire \efabless_subsystem.config_regs_i._2001_ ;
 wire \efabless_subsystem.config_regs_i._2002_ ;
 wire \efabless_subsystem.config_regs_i._2003_ ;
 wire \efabless_subsystem.config_regs_i._2004_ ;
 wire \efabless_subsystem.config_regs_i._2005_ ;
 wire \efabless_subsystem.config_regs_i._2006_ ;
 wire \efabless_subsystem.config_regs_i._2007_ ;
 wire \efabless_subsystem.config_regs_i._2008_ ;
 wire \efabless_subsystem.config_regs_i._2009_ ;
 wire \efabless_subsystem.config_regs_i._2010_ ;
 wire \efabless_subsystem.config_regs_i._2011_ ;
 wire \efabless_subsystem.config_regs_i._2012_ ;
 wire \efabless_subsystem.config_regs_i._2013_ ;
 wire \efabless_subsystem.config_regs_i._2014_ ;
 wire \efabless_subsystem.config_regs_i._2015_ ;
 wire \efabless_subsystem.config_regs_i._2046_ ;
 wire \efabless_subsystem.config_regs_i._2047_ ;
 wire \efabless_subsystem.config_regs_i._2048_ ;
 wire \efabless_subsystem.config_regs_i._2079_ ;
 wire \efabless_subsystem.config_regs_i._2080_ ;
 wire \efabless_subsystem.config_regs_i._2081_ ;
 wire \efabless_subsystem.config_regs_i._2088_ ;
 wire \efabless_subsystem.config_regs_i._2089_ ;
 wire \efabless_subsystem.config_regs_i._2090_ ;
 wire \efabless_subsystem.config_regs_i._2091_ ;
 wire \efabless_subsystem.config_regs_i._2092_ ;
 wire \efabless_subsystem.config_regs_i._2093_ ;
 wire \efabless_subsystem.config_regs_i._2094_ ;
 wire \efabless_subsystem.config_regs_i._2095_ ;
 wire \efabless_subsystem.config_regs_i._2096_ ;
 wire \efabless_subsystem.config_regs_i._2097_ ;
 wire \efabless_subsystem.config_regs_i._2098_ ;
 wire \efabless_subsystem.config_regs_i._2099_ ;
 wire \efabless_subsystem.config_regs_i._2100_ ;
 wire \efabless_subsystem.config_regs_i._2101_ ;
 wire \efabless_subsystem.config_regs_i._2102_ ;
 wire \efabless_subsystem.config_regs_i._2103_ ;
 wire \efabless_subsystem.config_regs_i._2104_ ;
 wire \efabless_subsystem.config_regs_i._2105_ ;
 wire \efabless_subsystem.config_regs_i._2109_ ;
 wire \efabless_subsystem.config_regs_i._2110_ ;
 wire \efabless_subsystem.config_regs_i._2111_ ;
 wire \efabless_subsystem.config_regs_i._2142_ ;
 wire \efabless_subsystem.config_regs_i._2143_ ;
 wire \efabless_subsystem.config_regs_i._2144_ ;
 wire \efabless_subsystem.config_regs_i._2175_ ;
 wire \efabless_subsystem.config_regs_i._2176_ ;
 wire \efabless_subsystem.config_regs_i._2177_ ;
 wire \efabless_subsystem.config_regs_i._2184_ ;
 wire \efabless_subsystem.config_regs_i._2185_ ;
 wire \efabless_subsystem.config_regs_i._2186_ ;
 wire \efabless_subsystem.config_regs_i._2187_ ;
 wire \efabless_subsystem.config_regs_i._2188_ ;
 wire \efabless_subsystem.config_regs_i._2189_ ;
 wire \efabless_subsystem.config_regs_i._2190_ ;
 wire \efabless_subsystem.config_regs_i._2191_ ;
 wire \efabless_subsystem.config_regs_i._2192_ ;
 wire \efabless_subsystem.config_regs_i._2193_ ;
 wire \efabless_subsystem.config_regs_i._2194_ ;
 wire \efabless_subsystem.config_regs_i._2195_ ;
 wire \efabless_subsystem.config_regs_i._2196_ ;
 wire \efabless_subsystem.config_regs_i._2197_ ;
 wire \efabless_subsystem.config_regs_i._2198_ ;
 wire \efabless_subsystem.config_regs_i._2199_ ;
 wire \efabless_subsystem.config_regs_i._2200_ ;
 wire \efabless_subsystem.config_regs_i._2201_ ;
 wire \efabless_subsystem.config_regs_i._2397_ ;
 wire \efabless_subsystem.config_regs_i._2398_ ;
 wire \efabless_subsystem.config_regs_i._2399_ ;
 wire \efabless_subsystem.config_regs_i._2400_ ;
 wire \efabless_subsystem.config_regs_i._2401_ ;
 wire \efabless_subsystem.config_regs_i._2402_ ;
 wire \efabless_subsystem.config_regs_i._2499_ ;
 wire \efabless_subsystem.config_regs_i._2500_ ;
 wire \efabless_subsystem.config_regs_i._2501_ ;
 wire \efabless_subsystem.config_regs_i._2502_ ;
 wire \efabless_subsystem.config_regs_i._2503_ ;
 wire \efabless_subsystem.config_regs_i._2504_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_d ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ;
 wire \efabless_subsystem.config_regs_i.count_enable_q_reg.srd ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[5] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[6] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._2_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424._1_ ;
 wire \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._01_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._02_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._03_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._05_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._06_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._07_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._08_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._09_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._10_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._11_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._12_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86._13_ ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[0] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[1] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[2] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[3] ;
 wire \efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[4] ;
 wire \efabless_subsystem.config_regs_i.done_ien_d ;
 wire \efabless_subsystem.config_regs_i.done_ien_q ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.done_ien_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_d ;
 wire \efabless_subsystem.config_regs_i.done_intr_q ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.done_intr_q_reg.srl ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg.d ;
 wire \efabless_subsystem.config_regs_i.global_ien_d ;
 wire \efabless_subsystem.config_regs_i.global_ien_q ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.global_ien_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.idle_d ;
 wire \efabless_subsystem.config_regs_i.idle_q ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg.srd ;
 wire \efabless_subsystem.config_regs_i.idle_q_reg.srl ;
 wire \efabless_subsystem.config_regs_i.mem_mode_d ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.mem_mode_q_reg.q ;
 wire \efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ;
 wire \efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_auto_restart_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_done_ien_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_global_ien_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_idle_d_379_18.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_mem_mode_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g29.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_rden_198_21.ctl ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.ctl[1] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_127.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_136.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_146.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_156.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_166.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_176.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_186.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_195.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_205.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_215.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_225.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_235.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_245.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_255.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_265.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_275.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_284.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_293.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_303.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_313.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_323.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_333.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_343.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_353.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_363.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_373.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_383.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_393.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_403.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_413.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_423.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_312_21.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_357_26.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_358_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_21.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_628.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_636.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_644.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_652.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_660.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_668.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_676.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_684.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_692.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_700.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_708.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_716.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_624.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_632.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_640.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_648.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_656.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_664.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_672.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_680.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_688.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_696.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_704.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_712.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_21.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_876.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_882.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_888.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_894.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_900.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_906.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_912.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_918.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_924.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_930.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_936.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_942.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_26.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_874.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_880.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_886.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_892.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_898.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_904.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_910.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_916.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_922.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_928.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_934.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_940.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_873.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_879.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_885.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_891.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_897.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_903.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_909.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_915.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_921.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_927.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_933.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_939.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1064.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1070.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1076.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1082.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1088.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1094.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1100.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1106.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_21.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1062.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1068.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1074.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1080.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1086.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1092.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1098.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1104.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_26.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1061.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1067.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1073.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1079.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1085.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1091.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1097.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1103.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.z ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1252.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1258.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1264.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1270.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1276.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1282.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1288.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1294.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_21.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1250.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1256.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1262.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1268.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1274.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1280.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1286.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1292.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_26.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1249.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1255.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1261.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1267.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1273.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1279.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1285.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1291.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1.z ;
 wire \efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_soft_rst_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_281_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.data0 ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.z ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_284_33.ctl ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_284_33.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_302_9.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_302_9.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_302_9.g1.z ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_306_17.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_306_17.g1.data1 ;
 wire \efabless_subsystem.config_regs_i.mux_start_d_312_21.ctl[0] ;
 wire \efabless_subsystem.config_regs_i.mux_wren_198_21.g1._0_ ;
 wire \efabless_subsystem.config_regs_i.o_doneintr ;
 wire \efabless_subsystem.config_regs_i.o_fifo_ptrs_set ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[0] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[10] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[11] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[12] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[1] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[2] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[3] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[4] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[5] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[6] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[7] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[8] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[9] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[0] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[10] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[11] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[12] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[1] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[2] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[3] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[4] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[5] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[6] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[7] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[8] ;
 wire \efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[9] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[0] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[1] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[2] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[3] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[4] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[5] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[6] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[7] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[8] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[0] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[1] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[2] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[3] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[4] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[5] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[6] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[7] ;
 wire \efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[8] ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.ready_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._06_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._00_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._01_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._02_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._03_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._04_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._05_ ;
 wire \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._06_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.soft_rst_q_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.start_q_prv_reg._06_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._00_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._01_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._02_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._03_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._04_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._05_ ;
 wire \efabless_subsystem.config_regs_i.start_q_reg._06_ ;
 wire \efabless_subsystem.core_stat_data_valid ;
 wire \efabless_subsystem.cpu_address[10] ;
 wire \efabless_subsystem.cpu_address[11] ;
 wire \efabless_subsystem.cpu_address[12] ;
 wire \efabless_subsystem.cpu_address[13] ;
 wire \efabless_subsystem.cpu_address[14] ;
 wire \efabless_subsystem.cpu_address[15] ;
 wire \efabless_subsystem.cpu_address[16] ;
 wire \efabless_subsystem.cpu_address[17] ;
 wire \efabless_subsystem.cpu_address[18] ;
 wire \efabless_subsystem.cpu_address[19] ;
 wire \efabless_subsystem.cpu_address[20] ;
 wire \efabless_subsystem.cpu_address[21] ;
 wire \efabless_subsystem.cpu_address[22] ;
 wire \efabless_subsystem.cpu_address[23] ;
 wire \efabless_subsystem.cpu_address[2] ;
 wire \efabless_subsystem.cpu_address[3] ;
 wire \efabless_subsystem.cpu_address[4] ;
 wire \efabless_subsystem.cpu_address[5] ;
 wire \efabless_subsystem.cpu_address[6] ;
 wire \efabless_subsystem.cpu_address[7] ;
 wire \efabless_subsystem.cpu_address[8] ;
 wire \efabless_subsystem.cpu_address[9] ;
 wire \efabless_subsystem.cpu_rden ;
 wire \efabless_subsystem.cpu_wdata[0] ;
 wire \efabless_subsystem.cpu_wdata[10] ;
 wire \efabless_subsystem.cpu_wdata[11] ;
 wire \efabless_subsystem.cpu_wdata[12] ;
 wire \efabless_subsystem.cpu_wdata[13] ;
 wire \efabless_subsystem.cpu_wdata[14] ;
 wire \efabless_subsystem.cpu_wdata[15] ;
 wire \efabless_subsystem.cpu_wdata[16] ;
 wire \efabless_subsystem.cpu_wdata[17] ;
 wire \efabless_subsystem.cpu_wdata[18] ;
 wire \efabless_subsystem.cpu_wdata[19] ;
 wire \efabless_subsystem.cpu_wdata[1] ;
 wire \efabless_subsystem.cpu_wdata[20] ;
 wire \efabless_subsystem.cpu_wdata[21] ;
 wire \efabless_subsystem.cpu_wdata[22] ;
 wire \efabless_subsystem.cpu_wdata[23] ;
 wire \efabless_subsystem.cpu_wdata[24] ;
 wire \efabless_subsystem.cpu_wdata[25] ;
 wire \efabless_subsystem.cpu_wdata[26] ;
 wire \efabless_subsystem.cpu_wdata[27] ;
 wire \efabless_subsystem.cpu_wdata[28] ;
 wire \efabless_subsystem.cpu_wdata[29] ;
 wire \efabless_subsystem.cpu_wdata[2] ;
 wire \efabless_subsystem.cpu_wdata[30] ;
 wire \efabless_subsystem.cpu_wdata[31] ;
 wire \efabless_subsystem.cpu_wdata[3] ;
 wire \efabless_subsystem.cpu_wdata[4] ;
 wire \efabless_subsystem.cpu_wdata[5] ;
 wire \efabless_subsystem.cpu_wdata[6] ;
 wire \efabless_subsystem.cpu_wdata[7] ;
 wire \efabless_subsystem.cpu_wdata[8] ;
 wire \efabless_subsystem.cpu_wdata[9] ;
 wire \efabless_subsystem.cpu_wmask[0] ;
 wire \efabless_subsystem.cpu_wmask[10] ;
 wire \efabless_subsystem.cpu_wmask[11] ;
 wire \efabless_subsystem.cpu_wmask[12] ;
 wire \efabless_subsystem.cpu_wmask[13] ;
 wire \efabless_subsystem.cpu_wmask[14] ;
 wire \efabless_subsystem.cpu_wmask[15] ;
 wire \efabless_subsystem.cpu_wmask[16] ;
 wire \efabless_subsystem.cpu_wmask[17] ;
 wire \efabless_subsystem.cpu_wmask[18] ;
 wire \efabless_subsystem.cpu_wmask[19] ;
 wire \efabless_subsystem.cpu_wmask[1] ;
 wire \efabless_subsystem.cpu_wmask[20] ;
 wire \efabless_subsystem.cpu_wmask[21] ;
 wire \efabless_subsystem.cpu_wmask[22] ;
 wire \efabless_subsystem.cpu_wmask[23] ;
 wire \efabless_subsystem.cpu_wmask[24] ;
 wire \efabless_subsystem.cpu_wmask[25] ;
 wire \efabless_subsystem.cpu_wmask[26] ;
 wire \efabless_subsystem.cpu_wmask[27] ;
 wire \efabless_subsystem.cpu_wmask[28] ;
 wire \efabless_subsystem.cpu_wmask[29] ;
 wire \efabless_subsystem.cpu_wmask[2] ;
 wire \efabless_subsystem.cpu_wmask[30] ;
 wire \efabless_subsystem.cpu_wmask[31] ;
 wire \efabless_subsystem.cpu_wmask[3] ;
 wire \efabless_subsystem.cpu_wmask[4] ;
 wire \efabless_subsystem.cpu_wmask[5] ;
 wire \efabless_subsystem.cpu_wmask[6] ;
 wire \efabless_subsystem.cpu_wmask[7] ;
 wire \efabless_subsystem.cpu_wmask[8] ;
 wire \efabless_subsystem.cpu_wmask[9] ;
 wire \efabless_subsystem.cpu_wren ;
 wire \efabless_subsystem.imem_acc_rdata_ready ;
 wire \efabless_subsystem.imem_acc_rdata_valid ;
 wire \efabless_subsystem.imem_address[0] ;
 wire \efabless_subsystem.imem_address[1] ;
 wire \efabless_subsystem.imem_address[2] ;
 wire \efabless_subsystem.imem_address[3] ;
 wire \efabless_subsystem.imem_address[4] ;
 wire \efabless_subsystem.imem_address[5] ;
 wire \efabless_subsystem.imem_rdata[0] ;
 wire \efabless_subsystem.imem_rdata[100] ;
 wire \efabless_subsystem.imem_rdata[101] ;
 wire \efabless_subsystem.imem_rdata[102] ;
 wire \efabless_subsystem.imem_rdata[103] ;
 wire \efabless_subsystem.imem_rdata[104] ;
 wire \efabless_subsystem.imem_rdata[105] ;
 wire \efabless_subsystem.imem_rdata[106] ;
 wire \efabless_subsystem.imem_rdata[107] ;
 wire \efabless_subsystem.imem_rdata[108] ;
 wire \efabless_subsystem.imem_rdata[109] ;
 wire \efabless_subsystem.imem_rdata[10] ;
 wire \efabless_subsystem.imem_rdata[110] ;
 wire \efabless_subsystem.imem_rdata[111] ;
 wire \efabless_subsystem.imem_rdata[112] ;
 wire \efabless_subsystem.imem_rdata[113] ;
 wire \efabless_subsystem.imem_rdata[114] ;
 wire \efabless_subsystem.imem_rdata[115] ;
 wire \efabless_subsystem.imem_rdata[116] ;
 wire \efabless_subsystem.imem_rdata[117] ;
 wire \efabless_subsystem.imem_rdata[118] ;
 wire \efabless_subsystem.imem_rdata[119] ;
 wire \efabless_subsystem.imem_rdata[11] ;
 wire \efabless_subsystem.imem_rdata[120] ;
 wire \efabless_subsystem.imem_rdata[121] ;
 wire \efabless_subsystem.imem_rdata[122] ;
 wire \efabless_subsystem.imem_rdata[123] ;
 wire \efabless_subsystem.imem_rdata[124] ;
 wire \efabless_subsystem.imem_rdata[125] ;
 wire \efabless_subsystem.imem_rdata[126] ;
 wire \efabless_subsystem.imem_rdata[127] ;
 wire \efabless_subsystem.imem_rdata[128] ;
 wire \efabless_subsystem.imem_rdata[129] ;
 wire \efabless_subsystem.imem_rdata[12] ;
 wire \efabless_subsystem.imem_rdata[130] ;
 wire \efabless_subsystem.imem_rdata[131] ;
 wire \efabless_subsystem.imem_rdata[132] ;
 wire \efabless_subsystem.imem_rdata[133] ;
 wire \efabless_subsystem.imem_rdata[134] ;
 wire \efabless_subsystem.imem_rdata[135] ;
 wire \efabless_subsystem.imem_rdata[136] ;
 wire \efabless_subsystem.imem_rdata[137] ;
 wire \efabless_subsystem.imem_rdata[138] ;
 wire \efabless_subsystem.imem_rdata[139] ;
 wire \efabless_subsystem.imem_rdata[13] ;
 wire \efabless_subsystem.imem_rdata[140] ;
 wire \efabless_subsystem.imem_rdata[141] ;
 wire \efabless_subsystem.imem_rdata[142] ;
 wire \efabless_subsystem.imem_rdata[143] ;
 wire \efabless_subsystem.imem_rdata[144] ;
 wire \efabless_subsystem.imem_rdata[145] ;
 wire \efabless_subsystem.imem_rdata[146] ;
 wire \efabless_subsystem.imem_rdata[147] ;
 wire \efabless_subsystem.imem_rdata[148] ;
 wire \efabless_subsystem.imem_rdata[149] ;
 wire \efabless_subsystem.imem_rdata[14] ;
 wire \efabless_subsystem.imem_rdata[150] ;
 wire \efabless_subsystem.imem_rdata[151] ;
 wire \efabless_subsystem.imem_rdata[152] ;
 wire \efabless_subsystem.imem_rdata[153] ;
 wire \efabless_subsystem.imem_rdata[154] ;
 wire \efabless_subsystem.imem_rdata[155] ;
 wire \efabless_subsystem.imem_rdata[156] ;
 wire \efabless_subsystem.imem_rdata[157] ;
 wire \efabless_subsystem.imem_rdata[158] ;
 wire \efabless_subsystem.imem_rdata[159] ;
 wire \efabless_subsystem.imem_rdata[15] ;
 wire \efabless_subsystem.imem_rdata[160] ;
 wire \efabless_subsystem.imem_rdata[161] ;
 wire \efabless_subsystem.imem_rdata[162] ;
 wire \efabless_subsystem.imem_rdata[163] ;
 wire \efabless_subsystem.imem_rdata[164] ;
 wire \efabless_subsystem.imem_rdata[165] ;
 wire \efabless_subsystem.imem_rdata[166] ;
 wire \efabless_subsystem.imem_rdata[167] ;
 wire \efabless_subsystem.imem_rdata[168] ;
 wire \efabless_subsystem.imem_rdata[169] ;
 wire \efabless_subsystem.imem_rdata[16] ;
 wire \efabless_subsystem.imem_rdata[170] ;
 wire \efabless_subsystem.imem_rdata[171] ;
 wire \efabless_subsystem.imem_rdata[172] ;
 wire \efabless_subsystem.imem_rdata[173] ;
 wire \efabless_subsystem.imem_rdata[174] ;
 wire \efabless_subsystem.imem_rdata[175] ;
 wire \efabless_subsystem.imem_rdata[176] ;
 wire \efabless_subsystem.imem_rdata[177] ;
 wire \efabless_subsystem.imem_rdata[178] ;
 wire \efabless_subsystem.imem_rdata[179] ;
 wire \efabless_subsystem.imem_rdata[17] ;
 wire \efabless_subsystem.imem_rdata[180] ;
 wire \efabless_subsystem.imem_rdata[181] ;
 wire \efabless_subsystem.imem_rdata[182] ;
 wire \efabless_subsystem.imem_rdata[183] ;
 wire \efabless_subsystem.imem_rdata[184] ;
 wire \efabless_subsystem.imem_rdata[185] ;
 wire \efabless_subsystem.imem_rdata[186] ;
 wire \efabless_subsystem.imem_rdata[187] ;
 wire \efabless_subsystem.imem_rdata[188] ;
 wire \efabless_subsystem.imem_rdata[189] ;
 wire \efabless_subsystem.imem_rdata[18] ;
 wire \efabless_subsystem.imem_rdata[190] ;
 wire \efabless_subsystem.imem_rdata[191] ;
 wire \efabless_subsystem.imem_rdata[192] ;
 wire \efabless_subsystem.imem_rdata[193] ;
 wire \efabless_subsystem.imem_rdata[194] ;
 wire \efabless_subsystem.imem_rdata[195] ;
 wire \efabless_subsystem.imem_rdata[196] ;
 wire \efabless_subsystem.imem_rdata[19] ;
 wire \efabless_subsystem.imem_rdata[1] ;
 wire \efabless_subsystem.imem_rdata[20] ;
 wire \efabless_subsystem.imem_rdata[21] ;
 wire \efabless_subsystem.imem_rdata[22] ;
 wire \efabless_subsystem.imem_rdata[23] ;
 wire \efabless_subsystem.imem_rdata[24] ;
 wire \efabless_subsystem.imem_rdata[25] ;
 wire \efabless_subsystem.imem_rdata[26] ;
 wire \efabless_subsystem.imem_rdata[27] ;
 wire \efabless_subsystem.imem_rdata[28] ;
 wire \efabless_subsystem.imem_rdata[29] ;
 wire \efabless_subsystem.imem_rdata[2] ;
 wire \efabless_subsystem.imem_rdata[30] ;
 wire \efabless_subsystem.imem_rdata[31] ;
 wire \efabless_subsystem.imem_rdata[32] ;
 wire \efabless_subsystem.imem_rdata[33] ;
 wire \efabless_subsystem.imem_rdata[34] ;
 wire \efabless_subsystem.imem_rdata[35] ;
 wire \efabless_subsystem.imem_rdata[36] ;
 wire \efabless_subsystem.imem_rdata[37] ;
 wire \efabless_subsystem.imem_rdata[38] ;
 wire \efabless_subsystem.imem_rdata[39] ;
 wire \efabless_subsystem.imem_rdata[3] ;
 wire \efabless_subsystem.imem_rdata[40] ;
 wire \efabless_subsystem.imem_rdata[41] ;
 wire \efabless_subsystem.imem_rdata[42] ;
 wire \efabless_subsystem.imem_rdata[43] ;
 wire \efabless_subsystem.imem_rdata[44] ;
 wire \efabless_subsystem.imem_rdata[45] ;
 wire \efabless_subsystem.imem_rdata[46] ;
 wire \efabless_subsystem.imem_rdata[47] ;
 wire \efabless_subsystem.imem_rdata[48] ;
 wire \efabless_subsystem.imem_rdata[49] ;
 wire \efabless_subsystem.imem_rdata[4] ;
 wire \efabless_subsystem.imem_rdata[50] ;
 wire \efabless_subsystem.imem_rdata[51] ;
 wire \efabless_subsystem.imem_rdata[52] ;
 wire \efabless_subsystem.imem_rdata[53] ;
 wire \efabless_subsystem.imem_rdata[54] ;
 wire \efabless_subsystem.imem_rdata[55] ;
 wire \efabless_subsystem.imem_rdata[56] ;
 wire \efabless_subsystem.imem_rdata[57] ;
 wire \efabless_subsystem.imem_rdata[58] ;
 wire \efabless_subsystem.imem_rdata[59] ;
 wire \efabless_subsystem.imem_rdata[5] ;
 wire \efabless_subsystem.imem_rdata[60] ;
 wire \efabless_subsystem.imem_rdata[61] ;
 wire \efabless_subsystem.imem_rdata[62] ;
 wire \efabless_subsystem.imem_rdata[63] ;
 wire \efabless_subsystem.imem_rdata[64] ;
 wire \efabless_subsystem.imem_rdata[65] ;
 wire \efabless_subsystem.imem_rdata[66] ;
 wire \efabless_subsystem.imem_rdata[67] ;
 wire \efabless_subsystem.imem_rdata[68] ;
 wire \efabless_subsystem.imem_rdata[69] ;
 wire \efabless_subsystem.imem_rdata[6] ;
 wire \efabless_subsystem.imem_rdata[70] ;
 wire \efabless_subsystem.imem_rdata[71] ;
 wire \efabless_subsystem.imem_rdata[72] ;
 wire \efabless_subsystem.imem_rdata[73] ;
 wire \efabless_subsystem.imem_rdata[74] ;
 wire \efabless_subsystem.imem_rdata[75] ;
 wire \efabless_subsystem.imem_rdata[76] ;
 wire \efabless_subsystem.imem_rdata[77] ;
 wire \efabless_subsystem.imem_rdata[78] ;
 wire \efabless_subsystem.imem_rdata[79] ;
 wire \efabless_subsystem.imem_rdata[7] ;
 wire \efabless_subsystem.imem_rdata[80] ;
 wire \efabless_subsystem.imem_rdata[81] ;
 wire \efabless_subsystem.imem_rdata[82] ;
 wire \efabless_subsystem.imem_rdata[83] ;
 wire \efabless_subsystem.imem_rdata[84] ;
 wire \efabless_subsystem.imem_rdata[85] ;
 wire \efabless_subsystem.imem_rdata[86] ;
 wire \efabless_subsystem.imem_rdata[87] ;
 wire \efabless_subsystem.imem_rdata[88] ;
 wire \efabless_subsystem.imem_rdata[89] ;
 wire \efabless_subsystem.imem_rdata[8] ;
 wire \efabless_subsystem.imem_rdata[90] ;
 wire \efabless_subsystem.imem_rdata[91] ;
 wire \efabless_subsystem.imem_rdata[92] ;
 wire \efabless_subsystem.imem_rdata[93] ;
 wire \efabless_subsystem.imem_rdata[94] ;
 wire \efabless_subsystem.imem_rdata[95] ;
 wire \efabless_subsystem.imem_rdata[96] ;
 wire \efabless_subsystem.imem_rdata[97] ;
 wire \efabless_subsystem.imem_rdata[98] ;
 wire \efabless_subsystem.imem_rdata[99] ;
 wire \efabless_subsystem.imem_rdata[9] ;
 wire \efabless_subsystem.imem_rden ;
 wire \efabless_subsystem.imem_wdata[0] ;
 wire \efabless_subsystem.imem_wdata[100] ;
 wire \efabless_subsystem.imem_wdata[101] ;
 wire \efabless_subsystem.imem_wdata[102] ;
 wire \efabless_subsystem.imem_wdata[103] ;
 wire \efabless_subsystem.imem_wdata[104] ;
 wire \efabless_subsystem.imem_wdata[105] ;
 wire \efabless_subsystem.imem_wdata[106] ;
 wire \efabless_subsystem.imem_wdata[107] ;
 wire \efabless_subsystem.imem_wdata[108] ;
 wire \efabless_subsystem.imem_wdata[109] ;
 wire \efabless_subsystem.imem_wdata[10] ;
 wire \efabless_subsystem.imem_wdata[110] ;
 wire \efabless_subsystem.imem_wdata[111] ;
 wire \efabless_subsystem.imem_wdata[112] ;
 wire \efabless_subsystem.imem_wdata[113] ;
 wire \efabless_subsystem.imem_wdata[114] ;
 wire \efabless_subsystem.imem_wdata[115] ;
 wire \efabless_subsystem.imem_wdata[116] ;
 wire \efabless_subsystem.imem_wdata[117] ;
 wire \efabless_subsystem.imem_wdata[118] ;
 wire \efabless_subsystem.imem_wdata[119] ;
 wire \efabless_subsystem.imem_wdata[11] ;
 wire \efabless_subsystem.imem_wdata[120] ;
 wire \efabless_subsystem.imem_wdata[121] ;
 wire \efabless_subsystem.imem_wdata[122] ;
 wire \efabless_subsystem.imem_wdata[123] ;
 wire \efabless_subsystem.imem_wdata[124] ;
 wire \efabless_subsystem.imem_wdata[125] ;
 wire \efabless_subsystem.imem_wdata[126] ;
 wire \efabless_subsystem.imem_wdata[127] ;
 wire \efabless_subsystem.imem_wdata[128] ;
 wire \efabless_subsystem.imem_wdata[129] ;
 wire \efabless_subsystem.imem_wdata[12] ;
 wire \efabless_subsystem.imem_wdata[130] ;
 wire \efabless_subsystem.imem_wdata[131] ;
 wire \efabless_subsystem.imem_wdata[132] ;
 wire \efabless_subsystem.imem_wdata[133] ;
 wire \efabless_subsystem.imem_wdata[134] ;
 wire \efabless_subsystem.imem_wdata[135] ;
 wire \efabless_subsystem.imem_wdata[136] ;
 wire \efabless_subsystem.imem_wdata[137] ;
 wire \efabless_subsystem.imem_wdata[138] ;
 wire \efabless_subsystem.imem_wdata[139] ;
 wire \efabless_subsystem.imem_wdata[13] ;
 wire \efabless_subsystem.imem_wdata[140] ;
 wire \efabless_subsystem.imem_wdata[141] ;
 wire \efabless_subsystem.imem_wdata[142] ;
 wire \efabless_subsystem.imem_wdata[143] ;
 wire \efabless_subsystem.imem_wdata[144] ;
 wire \efabless_subsystem.imem_wdata[145] ;
 wire \efabless_subsystem.imem_wdata[146] ;
 wire \efabless_subsystem.imem_wdata[147] ;
 wire \efabless_subsystem.imem_wdata[148] ;
 wire \efabless_subsystem.imem_wdata[149] ;
 wire \efabless_subsystem.imem_wdata[14] ;
 wire \efabless_subsystem.imem_wdata[150] ;
 wire \efabless_subsystem.imem_wdata[151] ;
 wire \efabless_subsystem.imem_wdata[152] ;
 wire \efabless_subsystem.imem_wdata[153] ;
 wire \efabless_subsystem.imem_wdata[154] ;
 wire \efabless_subsystem.imem_wdata[155] ;
 wire \efabless_subsystem.imem_wdata[156] ;
 wire \efabless_subsystem.imem_wdata[157] ;
 wire \efabless_subsystem.imem_wdata[158] ;
 wire \efabless_subsystem.imem_wdata[159] ;
 wire \efabless_subsystem.imem_wdata[15] ;
 wire \efabless_subsystem.imem_wdata[160] ;
 wire \efabless_subsystem.imem_wdata[161] ;
 wire \efabless_subsystem.imem_wdata[162] ;
 wire \efabless_subsystem.imem_wdata[163] ;
 wire \efabless_subsystem.imem_wdata[164] ;
 wire \efabless_subsystem.imem_wdata[165] ;
 wire \efabless_subsystem.imem_wdata[166] ;
 wire \efabless_subsystem.imem_wdata[167] ;
 wire \efabless_subsystem.imem_wdata[168] ;
 wire \efabless_subsystem.imem_wdata[169] ;
 wire \efabless_subsystem.imem_wdata[16] ;
 wire \efabless_subsystem.imem_wdata[170] ;
 wire \efabless_subsystem.imem_wdata[171] ;
 wire \efabless_subsystem.imem_wdata[172] ;
 wire \efabless_subsystem.imem_wdata[173] ;
 wire \efabless_subsystem.imem_wdata[174] ;
 wire \efabless_subsystem.imem_wdata[175] ;
 wire \efabless_subsystem.imem_wdata[176] ;
 wire \efabless_subsystem.imem_wdata[177] ;
 wire \efabless_subsystem.imem_wdata[178] ;
 wire \efabless_subsystem.imem_wdata[179] ;
 wire \efabless_subsystem.imem_wdata[17] ;
 wire \efabless_subsystem.imem_wdata[180] ;
 wire \efabless_subsystem.imem_wdata[181] ;
 wire \efabless_subsystem.imem_wdata[182] ;
 wire \efabless_subsystem.imem_wdata[183] ;
 wire \efabless_subsystem.imem_wdata[184] ;
 wire \efabless_subsystem.imem_wdata[185] ;
 wire \efabless_subsystem.imem_wdata[186] ;
 wire \efabless_subsystem.imem_wdata[187] ;
 wire \efabless_subsystem.imem_wdata[188] ;
 wire \efabless_subsystem.imem_wdata[189] ;
 wire \efabless_subsystem.imem_wdata[18] ;
 wire \efabless_subsystem.imem_wdata[190] ;
 wire \efabless_subsystem.imem_wdata[191] ;
 wire \efabless_subsystem.imem_wdata[192] ;
 wire \efabless_subsystem.imem_wdata[193] ;
 wire \efabless_subsystem.imem_wdata[194] ;
 wire \efabless_subsystem.imem_wdata[195] ;
 wire \efabless_subsystem.imem_wdata[196] ;
 wire \efabless_subsystem.imem_wdata[19] ;
 wire \efabless_subsystem.imem_wdata[1] ;
 wire \efabless_subsystem.imem_wdata[20] ;
 wire \efabless_subsystem.imem_wdata[21] ;
 wire \efabless_subsystem.imem_wdata[22] ;
 wire \efabless_subsystem.imem_wdata[23] ;
 wire \efabless_subsystem.imem_wdata[24] ;
 wire \efabless_subsystem.imem_wdata[25] ;
 wire \efabless_subsystem.imem_wdata[26] ;
 wire \efabless_subsystem.imem_wdata[27] ;
 wire \efabless_subsystem.imem_wdata[28] ;
 wire \efabless_subsystem.imem_wdata[29] ;
 wire \efabless_subsystem.imem_wdata[2] ;
 wire \efabless_subsystem.imem_wdata[30] ;
 wire \efabless_subsystem.imem_wdata[31] ;
 wire \efabless_subsystem.imem_wdata[32] ;
 wire \efabless_subsystem.imem_wdata[33] ;
 wire \efabless_subsystem.imem_wdata[34] ;
 wire \efabless_subsystem.imem_wdata[35] ;
 wire \efabless_subsystem.imem_wdata[36] ;
 wire \efabless_subsystem.imem_wdata[37] ;
 wire \efabless_subsystem.imem_wdata[38] ;
 wire \efabless_subsystem.imem_wdata[39] ;
 wire \efabless_subsystem.imem_wdata[3] ;
 wire \efabless_subsystem.imem_wdata[40] ;
 wire \efabless_subsystem.imem_wdata[41] ;
 wire \efabless_subsystem.imem_wdata[42] ;
 wire \efabless_subsystem.imem_wdata[43] ;
 wire \efabless_subsystem.imem_wdata[44] ;
 wire \efabless_subsystem.imem_wdata[45] ;
 wire \efabless_subsystem.imem_wdata[46] ;
 wire \efabless_subsystem.imem_wdata[47] ;
 wire \efabless_subsystem.imem_wdata[48] ;
 wire \efabless_subsystem.imem_wdata[49] ;
 wire \efabless_subsystem.imem_wdata[4] ;
 wire \efabless_subsystem.imem_wdata[50] ;
 wire \efabless_subsystem.imem_wdata[51] ;
 wire \efabless_subsystem.imem_wdata[52] ;
 wire \efabless_subsystem.imem_wdata[53] ;
 wire \efabless_subsystem.imem_wdata[54] ;
 wire \efabless_subsystem.imem_wdata[55] ;
 wire \efabless_subsystem.imem_wdata[56] ;
 wire \efabless_subsystem.imem_wdata[57] ;
 wire \efabless_subsystem.imem_wdata[58] ;
 wire \efabless_subsystem.imem_wdata[59] ;
 wire \efabless_subsystem.imem_wdata[5] ;
 wire \efabless_subsystem.imem_wdata[60] ;
 wire \efabless_subsystem.imem_wdata[61] ;
 wire \efabless_subsystem.imem_wdata[62] ;
 wire \efabless_subsystem.imem_wdata[63] ;
 wire \efabless_subsystem.imem_wdata[64] ;
 wire \efabless_subsystem.imem_wdata[65] ;
 wire \efabless_subsystem.imem_wdata[66] ;
 wire \efabless_subsystem.imem_wdata[67] ;
 wire \efabless_subsystem.imem_wdata[68] ;
 wire \efabless_subsystem.imem_wdata[69] ;
 wire \efabless_subsystem.imem_wdata[6] ;
 wire \efabless_subsystem.imem_wdata[70] ;
 wire \efabless_subsystem.imem_wdata[71] ;
 wire \efabless_subsystem.imem_wdata[72] ;
 wire \efabless_subsystem.imem_wdata[73] ;
 wire \efabless_subsystem.imem_wdata[74] ;
 wire \efabless_subsystem.imem_wdata[75] ;
 wire \efabless_subsystem.imem_wdata[76] ;
 wire \efabless_subsystem.imem_wdata[77] ;
 wire \efabless_subsystem.imem_wdata[78] ;
 wire \efabless_subsystem.imem_wdata[79] ;
 wire \efabless_subsystem.imem_wdata[7] ;
 wire \efabless_subsystem.imem_wdata[80] ;
 wire \efabless_subsystem.imem_wdata[81] ;
 wire \efabless_subsystem.imem_wdata[82] ;
 wire \efabless_subsystem.imem_wdata[83] ;
 wire \efabless_subsystem.imem_wdata[84] ;
 wire \efabless_subsystem.imem_wdata[85] ;
 wire \efabless_subsystem.imem_wdata[86] ;
 wire \efabless_subsystem.imem_wdata[87] ;
 wire \efabless_subsystem.imem_wdata[88] ;
 wire \efabless_subsystem.imem_wdata[89] ;
 wire \efabless_subsystem.imem_wdata[8] ;
 wire \efabless_subsystem.imem_wdata[90] ;
 wire \efabless_subsystem.imem_wdata[91] ;
 wire \efabless_subsystem.imem_wdata[92] ;
 wire \efabless_subsystem.imem_wdata[93] ;
 wire \efabless_subsystem.imem_wdata[94] ;
 wire \efabless_subsystem.imem_wdata[95] ;
 wire \efabless_subsystem.imem_wdata[96] ;
 wire \efabless_subsystem.imem_wdata[97] ;
 wire \efabless_subsystem.imem_wdata[98] ;
 wire \efabless_subsystem.imem_wdata[99] ;
 wire \efabless_subsystem.imem_wdata[9] ;
 wire \efabless_subsystem.imem_wmask[0] ;
 wire \efabless_subsystem.imem_wmask[104] ;
 wire \efabless_subsystem.imem_wmask[112] ;
 wire \efabless_subsystem.imem_wmask[120] ;
 wire \efabless_subsystem.imem_wmask[128] ;
 wire \efabless_subsystem.imem_wmask[136] ;
 wire \efabless_subsystem.imem_wmask[144] ;
 wire \efabless_subsystem.imem_wmask[152] ;
 wire \efabless_subsystem.imem_wmask[160] ;
 wire \efabless_subsystem.imem_wmask[168] ;
 wire \efabless_subsystem.imem_wmask[16] ;
 wire \efabless_subsystem.imem_wmask[176] ;
 wire \efabless_subsystem.imem_wmask[184] ;
 wire \efabless_subsystem.imem_wmask[192] ;
 wire \efabless_subsystem.imem_wmask[24] ;
 wire \efabless_subsystem.imem_wmask[32] ;
 wire \efabless_subsystem.imem_wmask[40] ;
 wire \efabless_subsystem.imem_wmask[48] ;
 wire \efabless_subsystem.imem_wmask[56] ;
 wire \efabless_subsystem.imem_wmask[64] ;
 wire \efabless_subsystem.imem_wmask[72] ;
 wire \efabless_subsystem.imem_wmask[80] ;
 wire \efabless_subsystem.imem_wmask[88] ;
 wire \efabless_subsystem.imem_wmask[8] ;
 wire \efabless_subsystem.imem_wmask[96] ;
 wire \efabless_subsystem.imem_wren ;
 wire \efabless_subsystem.input_memory_i._000_ ;
 wire \efabless_subsystem.input_memory_i._001_ ;
 wire \efabless_subsystem.input_memory_i._002_ ;
 wire \efabless_subsystem.input_memory_i._003_ ;
 wire \efabless_subsystem.input_memory_i._004_ ;
 wire \efabless_subsystem.input_memory_i._005_ ;
 wire \efabless_subsystem.input_memory_i._006_ ;
 wire \efabless_subsystem.input_memory_i._007_ ;
 wire \efabless_subsystem.input_memory_i._008_ ;
 wire \efabless_subsystem.input_memory_i._009_ ;
 wire \efabless_subsystem.input_memory_i._010_ ;
 wire \efabless_subsystem.input_memory_i._011_ ;
 wire \efabless_subsystem.input_memory_i._012_ ;
 wire \efabless_subsystem.input_memory_i._013_ ;
 wire \efabless_subsystem.input_memory_i._014_ ;
 wire \efabless_subsystem.input_memory_i._015_ ;
 wire \efabless_subsystem.input_memory_i._016_ ;
 wire \efabless_subsystem.input_memory_i._017_ ;
 wire \efabless_subsystem.input_memory_i._018_ ;
 wire \efabless_subsystem.input_memory_i._019_ ;
 wire \efabless_subsystem.input_memory_i._020_ ;
 wire \efabless_subsystem.input_memory_i._021_ ;
 wire \efabless_subsystem.input_memory_i._022_ ;
 wire \efabless_subsystem.input_memory_i._023_ ;
 wire \efabless_subsystem.input_memory_i._024_ ;
 wire \efabless_subsystem.input_memory_i._025_ ;
 wire \efabless_subsystem.input_memory_i._026_ ;
 wire \efabless_subsystem.input_memory_i._027_ ;
 wire \efabless_subsystem.input_memory_i._028_ ;
 wire \efabless_subsystem.input_memory_i._029_ ;
 wire \efabless_subsystem.input_memory_i._030_ ;
 wire \efabless_subsystem.input_memory_i._031_ ;
 wire \efabless_subsystem.input_memory_i._032_ ;
 wire \efabless_subsystem.input_memory_i._033_ ;
 wire \efabless_subsystem.input_memory_i._034_ ;
 wire \efabless_subsystem.input_memory_i._035_ ;
 wire \efabless_subsystem.input_memory_i._036_ ;
 wire \efabless_subsystem.input_memory_i._037_ ;
 wire \efabless_subsystem.input_memory_i._038_ ;
 wire \efabless_subsystem.input_memory_i._039_ ;
 wire \efabless_subsystem.input_memory_i._040_ ;
 wire \efabless_subsystem.input_memory_i._041_ ;
 wire \efabless_subsystem.input_memory_i._042_ ;
 wire \efabless_subsystem.input_memory_i._043_ ;
 wire \efabless_subsystem.input_memory_i._044_ ;
 wire \efabless_subsystem.input_memory_i._045_ ;
 wire \efabless_subsystem.input_memory_i._046_ ;
 wire \efabless_subsystem.input_memory_i._047_ ;
 wire \efabless_subsystem.input_memory_i._048_ ;
 wire \efabless_subsystem.input_memory_i._049_ ;
 wire \efabless_subsystem.input_memory_i._050_ ;
 wire \efabless_subsystem.input_memory_i._051_ ;
 wire \efabless_subsystem.input_memory_i._052_ ;
 wire \efabless_subsystem.input_memory_i._053_ ;
 wire \efabless_subsystem.input_memory_i._054_ ;
 wire \efabless_subsystem.input_memory_i._055_ ;
 wire \efabless_subsystem.input_memory_i._056_ ;
 wire \efabless_subsystem.input_memory_i._057_ ;
 wire \efabless_subsystem.input_memory_i._058_ ;
 wire \efabless_subsystem.input_memory_i._059_ ;
 wire \efabless_subsystem.input_memory_i._060_ ;
 wire \efabless_subsystem.input_memory_i._061_ ;
 wire \efabless_subsystem.input_memory_i._062_ ;
 wire \efabless_subsystem.input_memory_i._063_ ;
 wire \efabless_subsystem.input_memory_i._064_ ;
 wire \efabless_subsystem.input_memory_i._065_ ;
 wire \efabless_subsystem.input_memory_i._066_ ;
 wire \efabless_subsystem.input_memory_i._067_ ;
 wire \efabless_subsystem.input_memory_i._068_ ;
 wire \efabless_subsystem.input_memory_i._069_ ;
 wire \efabless_subsystem.input_memory_i._070_ ;
 wire \efabless_subsystem.input_memory_i._071_ ;
 wire \efabless_subsystem.input_memory_i._072_ ;
 wire \efabless_subsystem.input_memory_i._073_ ;
 wire \efabless_subsystem.input_memory_i._074_ ;
 wire \efabless_subsystem.input_memory_i._075_ ;
 wire \efabless_subsystem.input_memory_i._076_ ;
 wire \efabless_subsystem.input_memory_i._077_ ;
 wire \efabless_subsystem.input_memory_i._078_ ;
 wire \efabless_subsystem.input_memory_i._079_ ;
 wire \efabless_subsystem.input_memory_i._080_ ;
 wire \efabless_subsystem.input_memory_i._081_ ;
 wire \efabless_subsystem.input_memory_i._082_ ;
 wire \efabless_subsystem.input_memory_i._083_ ;
 wire \efabless_subsystem.input_memory_i._084_ ;
 wire \efabless_subsystem.input_memory_i._085_ ;
 wire \efabless_subsystem.input_memory_i._086_ ;
 wire \efabless_subsystem.input_memory_i._087_ ;
 wire \efabless_subsystem.input_memory_i._088_ ;
 wire \efabless_subsystem.input_memory_i._089_ ;
 wire \efabless_subsystem.input_memory_i._090_ ;
 wire \efabless_subsystem.input_memory_i._091_ ;
 wire \efabless_subsystem.input_memory_i._092_ ;
 wire \efabless_subsystem.input_memory_i._093_ ;
 wire \efabless_subsystem.input_memory_i._094_ ;
 wire \efabless_subsystem.input_memory_i._095_ ;
 wire \efabless_subsystem.input_memory_i._096_ ;
 wire \efabless_subsystem.input_memory_i._097_ ;
 wire \efabless_subsystem.input_memory_i._098_ ;
 wire \efabless_subsystem.input_memory_i._099_ ;
 wire \efabless_subsystem.input_memory_i._100_ ;
 wire \efabless_subsystem.input_memory_i._101_ ;
 wire \efabless_subsystem.input_memory_i._102_ ;
 wire \efabless_subsystem.input_memory_i._103_ ;
 wire \efabless_subsystem.input_memory_i._104_ ;
 wire \efabless_subsystem.input_memory_i._105_ ;
 wire \efabless_subsystem.input_memory_i._106_ ;
 wire \efabless_subsystem.input_memory_i._107_ ;
 wire \efabless_subsystem.input_memory_i._108_ ;
 wire \efabless_subsystem.input_memory_i._109_ ;
 wire \efabless_subsystem.input_memory_i._110_ ;
 wire \efabless_subsystem.input_memory_i._111_ ;
 wire \efabless_subsystem.input_memory_i._112_ ;
 wire \efabless_subsystem.input_memory_i._113_ ;
 wire \efabless_subsystem.input_memory_i._114_ ;
 wire \efabless_subsystem.input_memory_i._115_ ;
 wire \efabless_subsystem.input_memory_i._116_ ;
 wire \efabless_subsystem.input_memory_i._117_ ;
 wire \efabless_subsystem.input_memory_i._118_ ;
 wire \efabless_subsystem.input_memory_i._119_ ;
 wire \efabless_subsystem.input_memory_i._120_ ;
 wire \efabless_subsystem.input_memory_i._121_ ;
 wire \efabless_subsystem.input_memory_i._122_ ;
 wire \efabless_subsystem.input_memory_i._123_ ;
 wire \efabless_subsystem.input_memory_i._124_ ;
 wire \efabless_subsystem.input_memory_i._125_ ;
 wire \efabless_subsystem.input_memory_i._126_ ;
 wire \efabless_subsystem.input_memory_i._127_ ;
 wire \efabless_subsystem.input_memory_i._128_ ;
 wire \efabless_subsystem.input_memory_i._129_ ;
 wire \efabless_subsystem.input_memory_i._130_ ;
 wire \efabless_subsystem.input_memory_i._131_ ;
 wire \efabless_subsystem.input_memory_i._132_ ;
 wire \efabless_subsystem.input_memory_i._133_ ;
 wire \efabless_subsystem.input_memory_i._134_ ;
 wire \efabless_subsystem.input_memory_i._135_ ;
 wire \efabless_subsystem.input_memory_i._136_ ;
 wire \efabless_subsystem.input_memory_i._137_ ;
 wire \efabless_subsystem.input_memory_i._138_ ;
 wire \efabless_subsystem.input_memory_i._139_ ;
 wire \efabless_subsystem.input_memory_i._140_ ;
 wire \efabless_subsystem.input_memory_i._141_ ;
 wire \efabless_subsystem.input_memory_i._142_ ;
 wire \efabless_subsystem.input_memory_i._143_ ;
 wire \efabless_subsystem.input_memory_i._144_ ;
 wire \efabless_subsystem.input_memory_i._145_ ;
 wire \efabless_subsystem.input_memory_i._146_ ;
 wire \efabless_subsystem.input_memory_i._147_ ;
 wire \efabless_subsystem.input_memory_i._148_ ;
 wire \efabless_subsystem.input_memory_i._149_ ;
 wire \efabless_subsystem.input_memory_i._150_ ;
 wire \efabless_subsystem.input_memory_i._151_ ;
 wire \efabless_subsystem.input_memory_i._152_ ;
 wire \efabless_subsystem.input_memory_i._153_ ;
 wire \efabless_subsystem.input_memory_i._154_ ;
 wire \efabless_subsystem.input_memory_i._155_ ;
 wire \efabless_subsystem.input_memory_i._156_ ;
 wire \efabless_subsystem.input_memory_i._157_ ;
 wire \efabless_subsystem.input_memory_i._158_ ;
 wire \efabless_subsystem.input_memory_i._159_ ;
 wire \efabless_subsystem.input_memory_i._160_ ;
 wire \efabless_subsystem.input_memory_i._161_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[0] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[10] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[11] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[12] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[1] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[2] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[3] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[4] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[5] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[6] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[7] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[8] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.A[9] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[0] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[10] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[11] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[12] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[1] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[2] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[3] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[4] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[5] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[6] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[7] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[8] ;
 wire \efabless_subsystem.input_memory_i.add_144_39.Z[9] ;
 wire \efabless_subsystem.input_memory_i.add_144_39._00_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._01_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._02_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._03_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._04_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._05_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._06_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._07_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._08_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._09_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._10_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._11_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._12_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._13_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._14_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._15_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._16_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._17_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._18_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._19_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._20_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._21_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._22_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._23_ ;
 wire \efabless_subsystem.input_memory_i.add_144_39._24_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[0] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[10] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[11] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[12] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[1] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[2] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[3] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[4] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[5] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[6] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[7] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[8] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.A[9] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[0] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[10] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[11] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[12] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[1] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[2] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[3] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[4] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[5] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[6] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[7] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[8] ;
 wire \efabless_subsystem.input_memory_i.add_149_37.Z[9] ;
 wire \efabless_subsystem.input_memory_i.add_149_37._00_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._01_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._02_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._03_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._04_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._05_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._06_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._07_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._08_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._09_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._10_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._11_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._12_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._13_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._14_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._15_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._16_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._17_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._18_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._19_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._20_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._21_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._22_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._23_ ;
 wire \efabless_subsystem.input_memory_i.add_149_37._24_ ;
 wire \efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[0] ;
 wire \efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[1] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[0] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[10] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[11] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[12] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[1] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[2] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[3] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[4] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[5] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[6] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[7] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[8] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.A[9] ;
 wire \efabless_subsystem.input_memory_i.eq_159_52.Z ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._00_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._01_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._02_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._03_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._04_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._05_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._06_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._07_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._08_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._09_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._10_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._11_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._12_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._13_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._14_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._15_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._16_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._17_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._18_ ;
 wire \efabless_subsystem.input_memory_i.eq_159_52._19_ ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[0] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[10] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[11] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[12] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[1] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[2] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[3] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[4] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[5] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[6] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[7] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[8] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.A[9] ;
 wire \efabless_subsystem.input_memory_i.eq_160_52.Z ;
 wire \efabless_subsystem.input_memory_i.eq_160_52._0_ ;
 wire \efabless_subsystem.input_memory_i.eq_160_52._1_ ;
 wire \efabless_subsystem.input_memory_i.eq_160_52._2_ ;
 wire \efabless_subsystem.input_memory_i.eq_160_52._3_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._00_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._01_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._02_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._03_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._04_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._05_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0]._06_ ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0].d ;
 wire \efabless_subsystem.input_memory_i.fifo_state_reg[0].sena ;
 wire \efabless_subsystem.input_memory_i.memory_addr[0] ;
 wire \efabless_subsystem.input_memory_i.memory_addr[1] ;
 wire \efabless_subsystem.input_memory_i.memory_addr[2] ;
 wire \efabless_subsystem.input_memory_i.memory_addr[3] ;
 wire \efabless_subsystem.input_memory_i.memory_addr[4] ;
 wire \efabless_subsystem.input_memory_i.memory_addr[5] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[0] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[100] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[101] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[102] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[103] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[104] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[105] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[106] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[107] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[108] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[109] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[10] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[110] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[111] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[112] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[113] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[114] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[115] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[116] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[117] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[118] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[119] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[11] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[120] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[121] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[122] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[123] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[124] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[125] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[126] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[127] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[128] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[129] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[12] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[130] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[131] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[132] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[133] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[134] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[135] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[136] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[137] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[138] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[139] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[13] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[140] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[141] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[142] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[143] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[144] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[145] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[146] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[147] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[148] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[149] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[14] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[150] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[151] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[152] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[153] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[154] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[155] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[156] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[157] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[158] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[159] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[15] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[160] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[161] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[162] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[163] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[164] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[165] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[166] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[167] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[168] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[169] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[16] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[170] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[171] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[172] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[173] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[174] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[175] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[176] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[177] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[178] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[179] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[17] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[180] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[181] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[182] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[183] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[184] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[185] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[186] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[187] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[188] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[189] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[18] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[190] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[191] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[192] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[193] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[194] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[195] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[196] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[19] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[1] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[20] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[21] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[22] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[23] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[24] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[25] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[26] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[27] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[28] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[29] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[2] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[30] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[31] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[32] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[33] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[34] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[35] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[36] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[37] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[38] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[39] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[3] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[40] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[41] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[42] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[43] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[44] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[45] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[46] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[47] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[48] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[49] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[4] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[50] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[51] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[52] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[53] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[54] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[55] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[56] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[57] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[58] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[59] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[5] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[60] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[61] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[62] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[63] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[64] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[65] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[66] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[67] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[68] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[69] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[6] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[70] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[71] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[72] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[73] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[74] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[75] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[76] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[77] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[78] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[79] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[7] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[80] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[81] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[82] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[83] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[84] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[85] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[86] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[87] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[88] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[89] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[8] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[90] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[91] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[92] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[93] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[94] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[95] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[96] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[97] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[98] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[99] ;
 wire \efabless_subsystem.input_memory_i.memory_wdata[9] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[0] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[10] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[11] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[12] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[13] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[14] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[15] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[16] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[17] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[18] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[19] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[1] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[20] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[21] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[22] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[23] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[24] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[2] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[3] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[4] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[5] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[6] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[7] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[8] ;
 wire \efabless_subsystem.input_memory_i.memory_wmask[9] ;
 wire \efabless_subsystem.input_memory_i.memory_wren ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g100._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g101._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g102._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g103._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g104._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g105._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g106._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g107._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g108._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g109._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g110._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g111._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g112._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g113._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g114._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g115._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g116._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g117._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g118._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g119._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g120._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g121._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g122._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g123._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g124._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g125._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g126._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g127._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g128._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g129._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g13._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g130._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g131._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g132._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g133._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g134._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g135._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g136._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g137._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g138._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g139._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g14._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g140._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g141._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g142._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g143._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g144._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g145._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g146._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g147._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g148._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g149._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g15._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g150._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g151._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g152._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g153._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g154._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g155._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g156._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g157._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g158._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g159._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g16._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g160._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g161._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g162._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g163._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g164._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g165._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g166._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g167._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g168._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g169._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g17._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g170._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g171._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g172._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g173._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g174._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g175._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g176._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g177._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g178._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g179._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g18._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g180._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g181._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g182._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g183._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g184._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g185._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g186._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g187._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g188._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g189._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g19._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g190._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g191._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g192._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g193._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g194._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g195._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g196._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g197._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g2._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g20._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g21._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g22._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g23._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g24._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g25._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g26._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g27._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g28._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g29._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g3._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g30._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g31._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g32._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g33._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g34._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g35._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g36._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g37._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g38._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g39._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g4._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g40._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g41._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g42._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g43._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g44._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g45._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g46._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g47._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g48._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g49._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g5._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g50._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g51._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g52._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g53._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g54._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g55._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g56._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g57._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g58._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g59._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g6._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g60._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g61._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g62._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g63._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g64._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g65._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g66._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g67._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g68._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g69._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g70._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g71._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g72._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g73._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g74._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g75._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g76._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g77._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g78._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g79._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g80._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g81._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g82._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g83._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g84._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g85._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g86._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g87._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g88._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g89._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g90._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g91._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g92._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g93._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g94._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g95._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g96._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g97._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g98._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_82_26.g99._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g13._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g14._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g15._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g16._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g17._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g18._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g19._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g2._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g20._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g21._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g22._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g23._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g24._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g25._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g3._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g4._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g5._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g6._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_83_26.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_84_26.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_84_26.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_84_26.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_84_26.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_84_26.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_84_26.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_85_26.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_85_26.g1.data1 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9.z ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g13._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g2._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g3._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g4._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g5._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g6._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9.data0 ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9.z ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g1._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g10._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g11._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g12._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g13._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g2._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g3._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g4._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g5._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g6._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g7._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g8._0_ ;
 wire \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g9._0_ ;
 wire \efabless_subsystem.input_memory_i.n_572 ;
 wire \efabless_subsystem.input_memory_i.n_573 ;
 wire \efabless_subsystem.input_memory_i.n_574 ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._06_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._00_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._01_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._02_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._03_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._04_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._05_ ;
 wire \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._06_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._00_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._01_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._02_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._03_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._04_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._05_ ;
 wire \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._06_ ;
 wire \efabless_subsystem.io_oeb ;
 wire \efabless_subsystem.io_out ;
 wire \efabless_subsystem.la_data_out[0] ;
 wire \efabless_subsystem.la_data_out[100] ;
 wire \efabless_subsystem.la_data_out[101] ;
 wire \efabless_subsystem.la_data_out[102] ;
 wire \efabless_subsystem.la_data_out[103] ;
 wire \efabless_subsystem.la_data_out[104] ;
 wire \efabless_subsystem.la_data_out[105] ;
 wire \efabless_subsystem.la_data_out[106] ;
 wire \efabless_subsystem.la_data_out[107] ;
 wire \efabless_subsystem.la_data_out[108] ;
 wire \efabless_subsystem.la_data_out[109] ;
 wire \efabless_subsystem.la_data_out[10] ;
 wire \efabless_subsystem.la_data_out[110] ;
 wire \efabless_subsystem.la_data_out[111] ;
 wire \efabless_subsystem.la_data_out[112] ;
 wire \efabless_subsystem.la_data_out[113] ;
 wire \efabless_subsystem.la_data_out[114] ;
 wire \efabless_subsystem.la_data_out[115] ;
 wire \efabless_subsystem.la_data_out[116] ;
 wire \efabless_subsystem.la_data_out[117] ;
 wire \efabless_subsystem.la_data_out[118] ;
 wire \efabless_subsystem.la_data_out[119] ;
 wire \efabless_subsystem.la_data_out[11] ;
 wire \efabless_subsystem.la_data_out[120] ;
 wire \efabless_subsystem.la_data_out[121] ;
 wire \efabless_subsystem.la_data_out[122] ;
 wire \efabless_subsystem.la_data_out[123] ;
 wire \efabless_subsystem.la_data_out[124] ;
 wire \efabless_subsystem.la_data_out[125] ;
 wire \efabless_subsystem.la_data_out[126] ;
 wire \efabless_subsystem.la_data_out[127] ;
 wire \efabless_subsystem.la_data_out[12] ;
 wire \efabless_subsystem.la_data_out[13] ;
 wire \efabless_subsystem.la_data_out[14] ;
 wire \efabless_subsystem.la_data_out[15] ;
 wire \efabless_subsystem.la_data_out[16] ;
 wire \efabless_subsystem.la_data_out[17] ;
 wire \efabless_subsystem.la_data_out[18] ;
 wire \efabless_subsystem.la_data_out[19] ;
 wire \efabless_subsystem.la_data_out[1] ;
 wire \efabless_subsystem.la_data_out[20] ;
 wire \efabless_subsystem.la_data_out[21] ;
 wire \efabless_subsystem.la_data_out[22] ;
 wire \efabless_subsystem.la_data_out[23] ;
 wire \efabless_subsystem.la_data_out[24] ;
 wire \efabless_subsystem.la_data_out[25] ;
 wire \efabless_subsystem.la_data_out[26] ;
 wire \efabless_subsystem.la_data_out[27] ;
 wire \efabless_subsystem.la_data_out[28] ;
 wire \efabless_subsystem.la_data_out[29] ;
 wire \efabless_subsystem.la_data_out[2] ;
 wire \efabless_subsystem.la_data_out[30] ;
 wire \efabless_subsystem.la_data_out[31] ;
 wire \efabless_subsystem.la_data_out[32] ;
 wire \efabless_subsystem.la_data_out[33] ;
 wire \efabless_subsystem.la_data_out[34] ;
 wire \efabless_subsystem.la_data_out[35] ;
 wire \efabless_subsystem.la_data_out[36] ;
 wire \efabless_subsystem.la_data_out[37] ;
 wire \efabless_subsystem.la_data_out[38] ;
 wire \efabless_subsystem.la_data_out[39] ;
 wire \efabless_subsystem.la_data_out[3] ;
 wire \efabless_subsystem.la_data_out[40] ;
 wire \efabless_subsystem.la_data_out[41] ;
 wire \efabless_subsystem.la_data_out[42] ;
 wire \efabless_subsystem.la_data_out[43] ;
 wire \efabless_subsystem.la_data_out[44] ;
 wire \efabless_subsystem.la_data_out[45] ;
 wire \efabless_subsystem.la_data_out[46] ;
 wire \efabless_subsystem.la_data_out[47] ;
 wire \efabless_subsystem.la_data_out[48] ;
 wire \efabless_subsystem.la_data_out[49] ;
 wire \efabless_subsystem.la_data_out[4] ;
 wire \efabless_subsystem.la_data_out[50] ;
 wire \efabless_subsystem.la_data_out[51] ;
 wire \efabless_subsystem.la_data_out[52] ;
 wire \efabless_subsystem.la_data_out[53] ;
 wire \efabless_subsystem.la_data_out[54] ;
 wire \efabless_subsystem.la_data_out[55] ;
 wire \efabless_subsystem.la_data_out[56] ;
 wire \efabless_subsystem.la_data_out[57] ;
 wire \efabless_subsystem.la_data_out[58] ;
 wire \efabless_subsystem.la_data_out[59] ;
 wire \efabless_subsystem.la_data_out[5] ;
 wire \efabless_subsystem.la_data_out[60] ;
 wire \efabless_subsystem.la_data_out[61] ;
 wire \efabless_subsystem.la_data_out[62] ;
 wire \efabless_subsystem.la_data_out[63] ;
 wire \efabless_subsystem.la_data_out[64] ;
 wire \efabless_subsystem.la_data_out[65] ;
 wire \efabless_subsystem.la_data_out[66] ;
 wire \efabless_subsystem.la_data_out[67] ;
 wire \efabless_subsystem.la_data_out[68] ;
 wire \efabless_subsystem.la_data_out[69] ;
 wire \efabless_subsystem.la_data_out[6] ;
 wire \efabless_subsystem.la_data_out[70] ;
 wire \efabless_subsystem.la_data_out[71] ;
 wire \efabless_subsystem.la_data_out[72] ;
 wire \efabless_subsystem.la_data_out[73] ;
 wire \efabless_subsystem.la_data_out[74] ;
 wire \efabless_subsystem.la_data_out[75] ;
 wire \efabless_subsystem.la_data_out[76] ;
 wire \efabless_subsystem.la_data_out[77] ;
 wire \efabless_subsystem.la_data_out[78] ;
 wire \efabless_subsystem.la_data_out[79] ;
 wire \efabless_subsystem.la_data_out[7] ;
 wire \efabless_subsystem.la_data_out[80] ;
 wire \efabless_subsystem.la_data_out[81] ;
 wire \efabless_subsystem.la_data_out[82] ;
 wire \efabless_subsystem.la_data_out[83] ;
 wire \efabless_subsystem.la_data_out[84] ;
 wire \efabless_subsystem.la_data_out[85] ;
 wire \efabless_subsystem.la_data_out[86] ;
 wire \efabless_subsystem.la_data_out[87] ;
 wire \efabless_subsystem.la_data_out[88] ;
 wire \efabless_subsystem.la_data_out[89] ;
 wire \efabless_subsystem.la_data_out[8] ;
 wire \efabless_subsystem.la_data_out[90] ;
 wire \efabless_subsystem.la_data_out[91] ;
 wire \efabless_subsystem.la_data_out[92] ;
 wire \efabless_subsystem.la_data_out[93] ;
 wire \efabless_subsystem.la_data_out[94] ;
 wire \efabless_subsystem.la_data_out[95] ;
 wire \efabless_subsystem.la_data_out[96] ;
 wire \efabless_subsystem.la_data_out[97] ;
 wire \efabless_subsystem.la_data_out[98] ;
 wire \efabless_subsystem.la_data_out[99] ;
 wire \efabless_subsystem.la_data_out[9] ;
 wire \efabless_subsystem.mmap_interconnect_i._0000_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0001_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0002_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0004_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0005_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0006_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0009_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0010_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0039_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0047_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0055_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0063_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0071_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0079_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0087_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0095_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0103_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0111_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0119_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0127_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0135_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0143_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0151_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0159_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0167_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0175_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0183_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0191_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0199_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0231_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0239_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0247_ ;
 wire \efabless_subsystem.mmap_interconnect_i._0255_ ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[0] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[10] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[11] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[12] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[13] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[14] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[15] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[16] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[17] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[18] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[19] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[1] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[20] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[21] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[2] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[3] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[4] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[5] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[6] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[7] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[8] ;
 wire \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[9] ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_105_36.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_105_36.g1._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_106_36.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_106_36.g1._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_107_36.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_107_36.g1._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_107_36.g1.z ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_111_36.g1._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_112_36.g1._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_112_36.g1.z ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g16._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g24._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g8._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g16._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g24._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g8._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g16._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g24._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g8._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g16._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g24._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g8._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g16._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g24._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g8._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.ctl ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g16._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g24._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g32._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g8._0_ ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_address[0] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_address[1] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_address[2] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_address[3] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_address[4] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[0] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[10] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[11] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[12] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[13] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[14] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[15] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[16] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[17] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[18] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[19] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[1] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[20] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[21] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[2] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[3] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[4] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[5] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[6] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[7] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[8] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[9] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[0] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[16] ;
 wire \efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[8] ;
 wire \efabless_subsystem.mux_276_38.g1._0_ ;
 wire \efabless_subsystem.mux_276_38.g1.data1 ;
 wire \efabless_subsystem.mux_277_38.g1._0_ ;
 wire \efabless_subsystem.o_irq[1] ;
 wire \efabless_subsystem.o_irq[2] ;
 wire \efabless_subsystem.reduction_memory_i._000_ ;
 wire \efabless_subsystem.reduction_memory_i._001_ ;
 wire \efabless_subsystem.reduction_memory_i._002_ ;
 wire \efabless_subsystem.reduction_memory_i._003_ ;
 wire \efabless_subsystem.reduction_memory_i._004_ ;
 wire \efabless_subsystem.reduction_memory_i._005_ ;
 wire \efabless_subsystem.reduction_memory_i._006_ ;
 wire \efabless_subsystem.reduction_memory_i._007_ ;
 wire \efabless_subsystem.reduction_memory_i._008_ ;
 wire \efabless_subsystem.reduction_memory_i._009_ ;
 wire \efabless_subsystem.reduction_memory_i._010_ ;
 wire \efabless_subsystem.reduction_memory_i._011_ ;
 wire \efabless_subsystem.reduction_memory_i._012_ ;
 wire \efabless_subsystem.reduction_memory_i._013_ ;
 wire \efabless_subsystem.reduction_memory_i._014_ ;
 wire \efabless_subsystem.reduction_memory_i._015_ ;
 wire \efabless_subsystem.reduction_memory_i._016_ ;
 wire \efabless_subsystem.reduction_memory_i._017_ ;
 wire \efabless_subsystem.reduction_memory_i._018_ ;
 wire \efabless_subsystem.reduction_memory_i._019_ ;
 wire \efabless_subsystem.reduction_memory_i._020_ ;
 wire \efabless_subsystem.reduction_memory_i._021_ ;
 wire \efabless_subsystem.reduction_memory_i._022_ ;
 wire \efabless_subsystem.reduction_memory_i._023_ ;
 wire \efabless_subsystem.reduction_memory_i._024_ ;
 wire \efabless_subsystem.reduction_memory_i._025_ ;
 wire \efabless_subsystem.reduction_memory_i._026_ ;
 wire \efabless_subsystem.reduction_memory_i._027_ ;
 wire \efabless_subsystem.reduction_memory_i._028_ ;
 wire \efabless_subsystem.reduction_memory_i._029_ ;
 wire \efabless_subsystem.reduction_memory_i._030_ ;
 wire \efabless_subsystem.reduction_memory_i._031_ ;
 wire \efabless_subsystem.reduction_memory_i._032_ ;
 wire \efabless_subsystem.reduction_memory_i._033_ ;
 wire \efabless_subsystem.reduction_memory_i._034_ ;
 wire \efabless_subsystem.reduction_memory_i._035_ ;
 wire \efabless_subsystem.reduction_memory_i._036_ ;
 wire \efabless_subsystem.reduction_memory_i._037_ ;
 wire \efabless_subsystem.reduction_memory_i._038_ ;
 wire \efabless_subsystem.reduction_memory_i._039_ ;
 wire \efabless_subsystem.reduction_memory_i._040_ ;
 wire \efabless_subsystem.reduction_memory_i._041_ ;
 wire \efabless_subsystem.reduction_memory_i._042_ ;
 wire \efabless_subsystem.reduction_memory_i._043_ ;
 wire \efabless_subsystem.reduction_memory_i._044_ ;
 wire \efabless_subsystem.reduction_memory_i._045_ ;
 wire \efabless_subsystem.reduction_memory_i._046_ ;
 wire \efabless_subsystem.reduction_memory_i._047_ ;
 wire \efabless_subsystem.reduction_memory_i._048_ ;
 wire \efabless_subsystem.reduction_memory_i._049_ ;
 wire \efabless_subsystem.reduction_memory_i._050_ ;
 wire \efabless_subsystem.reduction_memory_i._051_ ;
 wire \efabless_subsystem.reduction_memory_i._052_ ;
 wire \efabless_subsystem.reduction_memory_i._053_ ;
 wire \efabless_subsystem.reduction_memory_i._054_ ;
 wire \efabless_subsystem.reduction_memory_i._055_ ;
 wire \efabless_subsystem.reduction_memory_i._056_ ;
 wire \efabless_subsystem.reduction_memory_i._057_ ;
 wire \efabless_subsystem.reduction_memory_i._058_ ;
 wire \efabless_subsystem.reduction_memory_i._059_ ;
 wire \efabless_subsystem.reduction_memory_i._060_ ;
 wire \efabless_subsystem.reduction_memory_i._061_ ;
 wire \efabless_subsystem.reduction_memory_i._062_ ;
 wire \efabless_subsystem.reduction_memory_i._063_ ;
 wire \efabless_subsystem.reduction_memory_i._064_ ;
 wire \efabless_subsystem.reduction_memory_i._065_ ;
 wire \efabless_subsystem.reduction_memory_i._066_ ;
 wire \efabless_subsystem.reduction_memory_i._067_ ;
 wire \efabless_subsystem.reduction_memory_i._068_ ;
 wire \efabless_subsystem.reduction_memory_i._069_ ;
 wire \efabless_subsystem.reduction_memory_i._070_ ;
 wire \efabless_subsystem.reduction_memory_i._071_ ;
 wire \efabless_subsystem.reduction_memory_i._072_ ;
 wire \efabless_subsystem.reduction_memory_i._073_ ;
 wire \efabless_subsystem.reduction_memory_i._074_ ;
 wire \efabless_subsystem.reduction_memory_i._075_ ;
 wire \efabless_subsystem.reduction_memory_i._076_ ;
 wire \efabless_subsystem.reduction_memory_i._077_ ;
 wire \efabless_subsystem.reduction_memory_i._078_ ;
 wire \efabless_subsystem.reduction_memory_i._079_ ;
 wire \efabless_subsystem.reduction_memory_i._080_ ;
 wire \efabless_subsystem.reduction_memory_i._081_ ;
 wire \efabless_subsystem.reduction_memory_i._082_ ;
 wire \efabless_subsystem.reduction_memory_i._083_ ;
 wire \efabless_subsystem.reduction_memory_i._084_ ;
 wire \efabless_subsystem.reduction_memory_i._085_ ;
 wire \efabless_subsystem.reduction_memory_i._086_ ;
 wire \efabless_subsystem.reduction_memory_i._087_ ;
 wire \efabless_subsystem.reduction_memory_i._088_ ;
 wire \efabless_subsystem.reduction_memory_i._089_ ;
 wire \efabless_subsystem.reduction_memory_i._090_ ;
 wire \efabless_subsystem.reduction_memory_i._091_ ;
 wire \efabless_subsystem.reduction_memory_i._092_ ;
 wire \efabless_subsystem.reduction_memory_i._093_ ;
 wire \efabless_subsystem.reduction_memory_i._094_ ;
 wire \efabless_subsystem.reduction_memory_i._095_ ;
 wire \efabless_subsystem.reduction_memory_i._096_ ;
 wire \efabless_subsystem.reduction_memory_i._097_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[0] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[1] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[2] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[3] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[4] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[5] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[6] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[7] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.A[8] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[0] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[1] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[2] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[3] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[4] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[5] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[6] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[7] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39.Z[8] ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._00_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._01_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._02_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._03_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._04_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._05_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._06_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._07_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._08_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._09_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._10_ ;
 wire \efabless_subsystem.reduction_memory_i.add_144_39._11_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[0] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[1] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[2] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[3] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[4] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[5] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[6] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[7] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.A[8] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[0] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[1] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[2] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[3] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[4] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[5] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[6] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[7] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37.Z[8] ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._00_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._01_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._02_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._03_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._04_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._05_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._06_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._07_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._08_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._09_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._10_ ;
 wire \efabless_subsystem.reduction_memory_i.add_149_37._11_ ;
 wire \efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.in_0 ;
 wire \efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[0] ;
 wire \efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[1] ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0].d ;
 wire \efabless_subsystem.reduction_memory_i.fifo_state_reg[0].sena ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[0] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[1] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[2] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[3] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[4] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[5] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[6] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[7] ;
 wire \efabless_subsystem.reduction_memory_i.g17.Z[8] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[0] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[1] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[2] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[3] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[4] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[5] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[6] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[7] ;
 wire \efabless_subsystem.reduction_memory_i.g18.Z[8] ;
 wire \efabless_subsystem.reduction_memory_i.memory_addr[0] ;
 wire \efabless_subsystem.reduction_memory_i.memory_addr[1] ;
 wire \efabless_subsystem.reduction_memory_i.memory_addr[2] ;
 wire \efabless_subsystem.reduction_memory_i.memory_addr[3] ;
 wire \efabless_subsystem.reduction_memory_i.memory_addr[4] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[0] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[10] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[11] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[12] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[13] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[14] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[15] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[16] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[17] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[18] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[19] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[1] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[20] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[21] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[2] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[3] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[4] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[5] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[6] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[7] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[8] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wdata[9] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wmask[0] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wmask[1] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wmask[2] ;
 wire \efabless_subsystem.reduction_memory_i.memory_wren ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g10._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g11._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g12._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g13._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g14._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g15._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g16._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g17._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g18._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g19._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g2._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g20._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g21._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g22._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g3._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g4._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g5._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g6._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g7._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g8._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_82_26.g9._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_83_26.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_83_26.g2._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_83_26.g3._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_84_26.g4._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_84_26.g5._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_84_26.g6._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_84_26.g7._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_84_26.g8._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_85_26.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_85_26.g1.data1 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g2._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g3._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g4._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g5._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g6._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g7._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g8._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g9._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9.data0 ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9.z ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g1._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g2._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g3._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g4._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g5._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g6._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g7._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g8._0_ ;
 wire \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g9._0_ ;
 wire \efabless_subsystem.reduction_memory_i.n_160 ;
 wire \efabless_subsystem.reduction_memory_i.n_161 ;
 wire \efabless_subsystem.reduction_memory_i.n_162 ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._06_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._00_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._01_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._02_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._03_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._04_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._05_ ;
 wire \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._06_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._000_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._001_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._002_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._003_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._004_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._005_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._006_ ;
 wire \efabless_subsystem.wishbone_2mmap_i._007_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.ack_delayed ;
 wire \efabless_subsystem.wishbone_2mmap_i.add_88_47.A ;
 wire \efabless_subsystem.wishbone_2mmap_i.add_88_47.Z ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._00_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._01_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._02_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._03_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._04_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._05_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._06_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0].aclr ;
 wire \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0].d ;
 wire \efabless_subsystem.wishbone_2mmap_i.mux_ack_delayed_83_27.g1._0_ ;
 wire \efabless_subsystem.wishbone_2mmap_i.mux_latency_cnt_d_87_17.g1._0_ ;

 sky130_fd_sc_hd__conb_1 _000_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[1]));
 sky130_fd_sc_hd__conb_1 _001_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[2]));
 sky130_fd_sc_hd__conb_1 _002_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[3]));
 sky130_fd_sc_hd__conb_1 _003_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[4]));
 sky130_fd_sc_hd__conb_1 _004_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[5]));
 sky130_fd_sc_hd__conb_1 _005_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[6]));
 sky130_fd_sc_hd__conb_1 _006_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[7]));
 sky130_fd_sc_hd__conb_1 _007_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[8]));
 sky130_fd_sc_hd__conb_1 _008_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[9]));
 sky130_fd_sc_hd__conb_1 _009_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[10]));
 sky130_fd_sc_hd__conb_1 _010_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[11]));
 sky130_fd_sc_hd__conb_1 _011_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[12]));
 sky130_fd_sc_hd__conb_1 _012_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[13]));
 sky130_fd_sc_hd__conb_1 _013_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[14]));
 sky130_fd_sc_hd__conb_1 _014_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[15]));
 sky130_fd_sc_hd__conb_1 _015_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[16]));
 sky130_fd_sc_hd__conb_1 _016_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[17]));
 sky130_fd_sc_hd__conb_1 _017_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[18]));
 sky130_fd_sc_hd__conb_1 _018_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[19]));
 sky130_fd_sc_hd__conb_1 _019_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[20]));
 sky130_fd_sc_hd__conb_1 _020_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[21]));
 sky130_fd_sc_hd__conb_1 _021_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[22]));
 sky130_fd_sc_hd__conb_1 _022_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[23]));
 sky130_fd_sc_hd__conb_1 _023_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[24]));
 sky130_fd_sc_hd__conb_1 _024_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[25]));
 sky130_fd_sc_hd__conb_1 _025_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[26]));
 sky130_fd_sc_hd__conb_1 _026_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[27]));
 sky130_fd_sc_hd__conb_1 _027_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[28]));
 sky130_fd_sc_hd__conb_1 _028_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[29]));
 sky130_fd_sc_hd__conb_1 _029_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[30]));
 sky130_fd_sc_hd__conb_1 _030_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[31]));
 sky130_fd_sc_hd__conb_1 _031_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[32]));
 sky130_fd_sc_hd__conb_1 _032_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[33]));
 sky130_fd_sc_hd__conb_1 _033_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[34]));
 sky130_fd_sc_hd__conb_1 _034_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[35]));
 sky130_fd_sc_hd__conb_1 _035_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[36]));
 sky130_fd_sc_hd__conb_1 _036_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_oeb[37]));
 sky130_fd_sc_hd__conb_1 _037_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[0]));
 sky130_fd_sc_hd__conb_1 _038_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[2]));
 sky130_fd_sc_hd__conb_1 _039_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[3]));
 sky130_fd_sc_hd__conb_1 _040_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[4]));
 sky130_fd_sc_hd__conb_1 _041_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[5]));
 sky130_fd_sc_hd__conb_1 _042_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[6]));
 sky130_fd_sc_hd__conb_1 _043_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[7]));
 sky130_fd_sc_hd__conb_1 _044_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[8]));
 sky130_fd_sc_hd__conb_1 _045_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[9]));
 sky130_fd_sc_hd__conb_1 _046_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[10]));
 sky130_fd_sc_hd__conb_1 _047_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[11]));
 sky130_fd_sc_hd__conb_1 _048_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[12]));
 sky130_fd_sc_hd__conb_1 _049_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[13]));
 sky130_fd_sc_hd__conb_1 _050_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[14]));
 sky130_fd_sc_hd__conb_1 _051_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[15]));
 sky130_fd_sc_hd__conb_1 _052_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[16]));
 sky130_fd_sc_hd__conb_1 _053_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[17]));
 sky130_fd_sc_hd__conb_1 _054_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[18]));
 sky130_fd_sc_hd__conb_1 _055_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[19]));
 sky130_fd_sc_hd__conb_1 _056_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[20]));
 sky130_fd_sc_hd__conb_1 _057_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[21]));
 sky130_fd_sc_hd__conb_1 _058_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[22]));
 sky130_fd_sc_hd__conb_1 _059_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[23]));
 sky130_fd_sc_hd__conb_1 _060_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[24]));
 sky130_fd_sc_hd__conb_1 _061_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[25]));
 sky130_fd_sc_hd__conb_1 _062_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[26]));
 sky130_fd_sc_hd__conb_1 _063_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[27]));
 sky130_fd_sc_hd__conb_1 _064_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[28]));
 sky130_fd_sc_hd__conb_1 _065_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[29]));
 sky130_fd_sc_hd__conb_1 _066_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[30]));
 sky130_fd_sc_hd__conb_1 _067_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[31]));
 sky130_fd_sc_hd__conb_1 _068_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[32]));
 sky130_fd_sc_hd__conb_1 _069_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[33]));
 sky130_fd_sc_hd__conb_1 _070_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[34]));
 sky130_fd_sc_hd__conb_1 _071_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[35]));
 sky130_fd_sc_hd__conb_1 _072_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[36]));
 sky130_fd_sc_hd__conb_1 _073_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(io_out[37]));
 sky130_fd_sc_hd__conb_1 _074_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[0]));
 sky130_fd_sc_hd__conb_1 _075_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[1]));
 sky130_fd_sc_hd__conb_1 _076_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[2]));
 sky130_fd_sc_hd__conb_1 _077_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[3]));
 sky130_fd_sc_hd__conb_1 _078_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[4]));
 sky130_fd_sc_hd__conb_1 _079_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[5]));
 sky130_fd_sc_hd__conb_1 _080_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[6]));
 sky130_fd_sc_hd__conb_1 _081_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[7]));
 sky130_fd_sc_hd__conb_1 _082_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[8]));
 sky130_fd_sc_hd__conb_1 _083_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[9]));
 sky130_fd_sc_hd__conb_1 _084_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[10]));
 sky130_fd_sc_hd__conb_1 _085_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[11]));
 sky130_fd_sc_hd__conb_1 _086_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[12]));
 sky130_fd_sc_hd__conb_1 _087_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[13]));
 sky130_fd_sc_hd__conb_1 _088_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[14]));
 sky130_fd_sc_hd__conb_1 _089_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[15]));
 sky130_fd_sc_hd__conb_1 _090_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[16]));
 sky130_fd_sc_hd__conb_1 _091_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[17]));
 sky130_fd_sc_hd__conb_1 _092_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[18]));
 sky130_fd_sc_hd__conb_1 _093_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[19]));
 sky130_fd_sc_hd__conb_1 _094_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[20]));
 sky130_fd_sc_hd__conb_1 _095_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[21]));
 sky130_fd_sc_hd__conb_1 _096_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[22]));
 sky130_fd_sc_hd__conb_1 _097_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[23]));
 sky130_fd_sc_hd__conb_1 _098_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[24]));
 sky130_fd_sc_hd__conb_1 _099_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[25]));
 sky130_fd_sc_hd__conb_1 _100_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[26]));
 sky130_fd_sc_hd__conb_1 _101_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[27]));
 sky130_fd_sc_hd__conb_1 _102_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[28]));
 sky130_fd_sc_hd__conb_1 _103_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[29]));
 sky130_fd_sc_hd__conb_1 _104_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[30]));
 sky130_fd_sc_hd__conb_1 _105_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_2 _106_ (.A(\efabless_subsystem.io_oeb ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_oeb[0]));
 sky130_fd_sc_hd__buf_2 _107_ (.A(\efabless_subsystem.io_out ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 _108_ (.A(\efabless_subsystem.la_data_out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[0]));
 sky130_fd_sc_hd__buf_2 _109_ (.A(\efabless_subsystem.la_data_out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__buf_2 _110_ (.A(\efabless_subsystem.la_data_out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__buf_2 _111_ (.A(\efabless_subsystem.la_data_out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[3]));
 sky130_fd_sc_hd__buf_2 _112_ (.A(\efabless_subsystem.la_data_out[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__buf_2 _113_ (.A(\efabless_subsystem.la_data_out[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__buf_2 _114_ (.A(\efabless_subsystem.la_data_out[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__buf_2 _115_ (.A(\efabless_subsystem.la_data_out[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__buf_2 _116_ (.A(\efabless_subsystem.la_data_out[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__buf_2 _117_ (.A(\efabless_subsystem.la_data_out[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__buf_2 _118_ (.A(\efabless_subsystem.la_data_out[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__buf_2 _119_ (.A(\efabless_subsystem.la_data_out[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__buf_2 _120_ (.A(\efabless_subsystem.la_data_out[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[12]));
 sky130_fd_sc_hd__buf_2 _121_ (.A(\efabless_subsystem.la_data_out[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[13]));
 sky130_fd_sc_hd__buf_2 _122_ (.A(\efabless_subsystem.la_data_out[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[14]));
 sky130_fd_sc_hd__buf_2 _123_ (.A(\efabless_subsystem.la_data_out[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[15]));
 sky130_fd_sc_hd__buf_2 _124_ (.A(\efabless_subsystem.la_data_out[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[16]));
 sky130_fd_sc_hd__buf_2 _125_ (.A(\efabless_subsystem.la_data_out[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[17]));
 sky130_fd_sc_hd__buf_2 _126_ (.A(\efabless_subsystem.la_data_out[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[18]));
 sky130_fd_sc_hd__buf_2 _127_ (.A(\efabless_subsystem.la_data_out[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[19]));
 sky130_fd_sc_hd__buf_2 _128_ (.A(\efabless_subsystem.la_data_out[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[20]));
 sky130_fd_sc_hd__buf_2 _129_ (.A(\efabless_subsystem.la_data_out[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[21]));
 sky130_fd_sc_hd__buf_2 _130_ (.A(\efabless_subsystem.la_data_out[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[22]));
 sky130_fd_sc_hd__buf_2 _131_ (.A(\efabless_subsystem.la_data_out[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[23]));
 sky130_fd_sc_hd__buf_2 _132_ (.A(\efabless_subsystem.la_data_out[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[24]));
 sky130_fd_sc_hd__buf_2 _133_ (.A(\efabless_subsystem.la_data_out[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[25]));
 sky130_fd_sc_hd__buf_2 _134_ (.A(\efabless_subsystem.la_data_out[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[26]));
 sky130_fd_sc_hd__buf_2 _135_ (.A(\efabless_subsystem.la_data_out[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[27]));
 sky130_fd_sc_hd__buf_2 _136_ (.A(\efabless_subsystem.la_data_out[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[28]));
 sky130_fd_sc_hd__buf_2 _137_ (.A(\efabless_subsystem.la_data_out[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[29]));
 sky130_fd_sc_hd__buf_2 _138_ (.A(\efabless_subsystem.la_data_out[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[30]));
 sky130_fd_sc_hd__buf_2 _139_ (.A(\efabless_subsystem.la_data_out[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[31]));
 sky130_fd_sc_hd__buf_2 _140_ (.A(\efabless_subsystem.la_data_out[32] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__buf_2 _141_ (.A(\efabless_subsystem.la_data_out[33] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__buf_2 _142_ (.A(\efabless_subsystem.la_data_out[34] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__buf_2 _143_ (.A(\efabless_subsystem.la_data_out[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__buf_2 _144_ (.A(\efabless_subsystem.la_data_out[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__buf_2 _145_ (.A(\efabless_subsystem.la_data_out[37] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__buf_2 _146_ (.A(\efabless_subsystem.la_data_out[38] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__buf_2 _147_ (.A(\efabless_subsystem.la_data_out[39] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__buf_2 _148_ (.A(\efabless_subsystem.la_data_out[40] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[40]));
 sky130_fd_sc_hd__buf_2 _149_ (.A(\efabless_subsystem.la_data_out[41] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[41]));
 sky130_fd_sc_hd__buf_2 _150_ (.A(\efabless_subsystem.la_data_out[42] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[42]));
 sky130_fd_sc_hd__buf_2 _151_ (.A(\efabless_subsystem.la_data_out[43] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[43]));
 sky130_fd_sc_hd__buf_2 _152_ (.A(\efabless_subsystem.la_data_out[44] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[44]));
 sky130_fd_sc_hd__buf_2 _153_ (.A(\efabless_subsystem.la_data_out[45] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[45]));
 sky130_fd_sc_hd__buf_2 _154_ (.A(\efabless_subsystem.la_data_out[46] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[46]));
 sky130_fd_sc_hd__buf_2 _155_ (.A(\efabless_subsystem.la_data_out[47] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[47]));
 sky130_fd_sc_hd__buf_2 _156_ (.A(\efabless_subsystem.la_data_out[48] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[48]));
 sky130_fd_sc_hd__buf_2 _157_ (.A(\efabless_subsystem.la_data_out[49] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[49]));
 sky130_fd_sc_hd__buf_2 _158_ (.A(\efabless_subsystem.la_data_out[50] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[50]));
 sky130_fd_sc_hd__buf_2 _159_ (.A(\efabless_subsystem.la_data_out[51] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[51]));
 sky130_fd_sc_hd__buf_2 _160_ (.A(\efabless_subsystem.la_data_out[52] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[52]));
 sky130_fd_sc_hd__buf_2 _161_ (.A(\efabless_subsystem.la_data_out[53] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[53]));
 sky130_fd_sc_hd__buf_2 _162_ (.A(\efabless_subsystem.la_data_out[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[54]));
 sky130_fd_sc_hd__buf_2 _163_ (.A(\efabless_subsystem.la_data_out[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[55]));
 sky130_fd_sc_hd__buf_2 _164_ (.A(\efabless_subsystem.la_data_out[56] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[56]));
 sky130_fd_sc_hd__buf_2 _165_ (.A(\efabless_subsystem.la_data_out[57] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[57]));
 sky130_fd_sc_hd__buf_2 _166_ (.A(\efabless_subsystem.la_data_out[58] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[58]));
 sky130_fd_sc_hd__buf_2 _167_ (.A(\efabless_subsystem.la_data_out[59] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[59]));
 sky130_fd_sc_hd__buf_2 _168_ (.A(\efabless_subsystem.la_data_out[60] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[60]));
 sky130_fd_sc_hd__buf_2 _169_ (.A(\efabless_subsystem.la_data_out[61] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[61]));
 sky130_fd_sc_hd__buf_2 _170_ (.A(\efabless_subsystem.la_data_out[62] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[62]));
 sky130_fd_sc_hd__buf_2 _171_ (.A(\efabless_subsystem.la_data_out[63] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[63]));
 sky130_fd_sc_hd__buf_2 _172_ (.A(\efabless_subsystem.la_data_out[64] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[64]));
 sky130_fd_sc_hd__buf_2 _173_ (.A(\efabless_subsystem.la_data_out[65] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[65]));
 sky130_fd_sc_hd__buf_2 _174_ (.A(\efabless_subsystem.la_data_out[66] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[66]));
 sky130_fd_sc_hd__buf_2 _175_ (.A(\efabless_subsystem.la_data_out[67] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[67]));
 sky130_fd_sc_hd__buf_2 _176_ (.A(\efabless_subsystem.la_data_out[68] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[68]));
 sky130_fd_sc_hd__buf_2 _177_ (.A(\efabless_subsystem.la_data_out[69] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[69]));
 sky130_fd_sc_hd__buf_2 _178_ (.A(\efabless_subsystem.la_data_out[70] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[70]));
 sky130_fd_sc_hd__buf_2 _179_ (.A(\efabless_subsystem.la_data_out[71] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[71]));
 sky130_fd_sc_hd__buf_2 _180_ (.A(\efabless_subsystem.la_data_out[72] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[72]));
 sky130_fd_sc_hd__buf_2 _181_ (.A(\efabless_subsystem.la_data_out[73] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[73]));
 sky130_fd_sc_hd__buf_2 _182_ (.A(\efabless_subsystem.la_data_out[74] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[74]));
 sky130_fd_sc_hd__buf_2 _183_ (.A(\efabless_subsystem.la_data_out[75] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[75]));
 sky130_fd_sc_hd__buf_2 _184_ (.A(\efabless_subsystem.la_data_out[76] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[76]));
 sky130_fd_sc_hd__buf_2 _185_ (.A(\efabless_subsystem.la_data_out[77] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[77]));
 sky130_fd_sc_hd__buf_2 _186_ (.A(\efabless_subsystem.la_data_out[78] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[78]));
 sky130_fd_sc_hd__buf_2 _187_ (.A(\efabless_subsystem.la_data_out[79] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[79]));
 sky130_fd_sc_hd__buf_2 _188_ (.A(\efabless_subsystem.la_data_out[80] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[80]));
 sky130_fd_sc_hd__buf_2 _189_ (.A(\efabless_subsystem.la_data_out[81] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[81]));
 sky130_fd_sc_hd__buf_2 _190_ (.A(\efabless_subsystem.la_data_out[82] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[82]));
 sky130_fd_sc_hd__buf_2 _191_ (.A(\efabless_subsystem.la_data_out[83] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[83]));
 sky130_fd_sc_hd__buf_2 _192_ (.A(\efabless_subsystem.la_data_out[84] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[84]));
 sky130_fd_sc_hd__buf_2 _193_ (.A(\efabless_subsystem.la_data_out[85] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[85]));
 sky130_fd_sc_hd__buf_2 _194_ (.A(\efabless_subsystem.la_data_out[86] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[86]));
 sky130_fd_sc_hd__buf_2 _195_ (.A(\efabless_subsystem.la_data_out[87] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[87]));
 sky130_fd_sc_hd__buf_2 _196_ (.A(\efabless_subsystem.la_data_out[88] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[88]));
 sky130_fd_sc_hd__buf_2 _197_ (.A(\efabless_subsystem.la_data_out[89] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[89]));
 sky130_fd_sc_hd__buf_2 _198_ (.A(\efabless_subsystem.la_data_out[90] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[90]));
 sky130_fd_sc_hd__buf_2 _199_ (.A(\efabless_subsystem.la_data_out[91] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[91]));
 sky130_fd_sc_hd__buf_2 _200_ (.A(\efabless_subsystem.la_data_out[92] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[92]));
 sky130_fd_sc_hd__buf_2 _201_ (.A(\efabless_subsystem.la_data_out[93] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[93]));
 sky130_fd_sc_hd__buf_2 _202_ (.A(\efabless_subsystem.la_data_out[94] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[94]));
 sky130_fd_sc_hd__buf_2 _203_ (.A(\efabless_subsystem.la_data_out[95] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[95]));
 sky130_fd_sc_hd__buf_2 _204_ (.A(\efabless_subsystem.la_data_out[96] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[96]));
 sky130_fd_sc_hd__buf_2 _205_ (.A(\efabless_subsystem.la_data_out[97] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[97]));
 sky130_fd_sc_hd__buf_2 _206_ (.A(\efabless_subsystem.la_data_out[98] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[98]));
 sky130_fd_sc_hd__buf_2 _207_ (.A(\efabless_subsystem.la_data_out[99] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[99]));
 sky130_fd_sc_hd__buf_2 _208_ (.A(\efabless_subsystem.la_data_out[100] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[100]));
 sky130_fd_sc_hd__buf_2 _209_ (.A(\efabless_subsystem.la_data_out[101] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[101]));
 sky130_fd_sc_hd__buf_2 _210_ (.A(\efabless_subsystem.la_data_out[102] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[102]));
 sky130_fd_sc_hd__buf_2 _211_ (.A(\efabless_subsystem.la_data_out[103] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[103]));
 sky130_fd_sc_hd__buf_2 _212_ (.A(\efabless_subsystem.la_data_out[104] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[104]));
 sky130_fd_sc_hd__buf_2 _213_ (.A(\efabless_subsystem.la_data_out[105] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[105]));
 sky130_fd_sc_hd__buf_2 _214_ (.A(\efabless_subsystem.la_data_out[106] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[106]));
 sky130_fd_sc_hd__buf_2 _215_ (.A(\efabless_subsystem.la_data_out[107] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[107]));
 sky130_fd_sc_hd__buf_2 _216_ (.A(\efabless_subsystem.la_data_out[108] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[108]));
 sky130_fd_sc_hd__buf_2 _217_ (.A(\efabless_subsystem.la_data_out[109] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[109]));
 sky130_fd_sc_hd__buf_2 _218_ (.A(\efabless_subsystem.la_data_out[110] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[110]));
 sky130_fd_sc_hd__buf_2 _219_ (.A(\efabless_subsystem.la_data_out[111] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[111]));
 sky130_fd_sc_hd__buf_2 _220_ (.A(\efabless_subsystem.la_data_out[112] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[112]));
 sky130_fd_sc_hd__buf_2 _221_ (.A(\efabless_subsystem.la_data_out[113] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[113]));
 sky130_fd_sc_hd__buf_2 _222_ (.A(\efabless_subsystem.la_data_out[114] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[114]));
 sky130_fd_sc_hd__buf_2 _223_ (.A(\efabless_subsystem.la_data_out[115] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[115]));
 sky130_fd_sc_hd__buf_2 _224_ (.A(\efabless_subsystem.la_data_out[116] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[116]));
 sky130_fd_sc_hd__buf_2 _225_ (.A(\efabless_subsystem.la_data_out[117] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[117]));
 sky130_fd_sc_hd__buf_2 _226_ (.A(\efabless_subsystem.la_data_out[118] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[118]));
 sky130_fd_sc_hd__buf_2 _227_ (.A(\efabless_subsystem.la_data_out[119] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[119]));
 sky130_fd_sc_hd__buf_2 _228_ (.A(\efabless_subsystem.la_data_out[120] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[120]));
 sky130_fd_sc_hd__buf_2 _229_ (.A(\efabless_subsystem.la_data_out[121] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[121]));
 sky130_fd_sc_hd__buf_2 _230_ (.A(\efabless_subsystem.la_data_out[122] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[122]));
 sky130_fd_sc_hd__buf_2 _231_ (.A(\efabless_subsystem.la_data_out[123] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[123]));
 sky130_fd_sc_hd__buf_2 _232_ (.A(\efabless_subsystem.la_data_out[124] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[124]));
 sky130_fd_sc_hd__buf_2 _233_ (.A(\efabless_subsystem.la_data_out[125] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[125]));
 sky130_fd_sc_hd__buf_2 _234_ (.A(\efabless_subsystem.la_data_out[126] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[126]));
 sky130_fd_sc_hd__buf_2 _235_ (.A(\efabless_subsystem.la_data_out[127] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(la_data_out[127]));
 sky130_fd_sc_hd__buf_2 _236_ (.A(\efabless_subsystem.config_regs_i.o_doneintr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(user_irq[0]));
 sky130_fd_sc_hd__buf_2 _237_ (.A(\efabless_subsystem.o_irq[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(user_irq[1]));
 sky130_fd_sc_hd__buf_2 _238_ (.A(\efabless_subsystem.o_irq[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(user_irq[2]));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem._224_  (.A(\efabless_subsystem.imem_acc_rdata_valid ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2.z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem._000_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem._225_  (.A(\efabless_subsystem._000_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.i_array_shftsgn_valid ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem._226_  (.A(\efabless_subsystem.imem_acc_rdata_valid ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2.z ),
    .C(\efabless_subsystem.core_stat_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem._001_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem._227_  (.A(\efabless_subsystem._001_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mux_276_38.g1.data1 ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem._228_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2.z ),
    .B(\efabless_subsystem.compute_core_i.ifmap_regs_i.o_ready ),
    .C(\efabless_subsystem.compute_core_i.o_weight_ready ),
    .D(\efabless_subsystem.compute_core_i.o_array_shftsgn_ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem._002_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem._229_  (.A(\efabless_subsystem._002_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_acc_rdata_ready ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._230_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._003_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._231_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._004_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._232_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._005_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._233_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._006_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._234_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._007_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._235_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._008_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._236_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._009_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._237_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._010_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._238_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._011_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._239_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._012_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._240_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._013_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._241_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._014_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._242_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._015_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._243_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._016_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._244_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._017_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._245_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._018_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._246_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._019_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._247_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._020_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._248_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._021_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._249_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._022_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._250_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._023_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._251_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._024_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._252_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._025_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._253_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._026_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._254_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._027_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._255_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._028_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._256_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._029_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._257_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._030_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._258_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._031_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._259_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._032_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._260_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._033_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._261_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._034_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._262_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._035_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._263_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._036_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._264_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._037_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._265_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._038_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._266_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._039_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._267_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._040_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._268_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._041_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._269_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._042_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._270_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._043_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._271_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._272_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._045_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._273_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._274_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._275_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._276_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._049_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._277_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._050_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._278_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._051_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._279_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._052_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._280_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._053_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._281_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._054_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._282_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._055_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._283_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._056_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._284_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._057_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._285_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._058_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._286_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._059_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._287_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._060_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._288_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._061_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._289_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._062_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._290_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._063_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._291_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._064_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._292_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._065_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._293_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._066_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._294_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._067_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._295_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._068_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._296_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._069_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._297_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._070_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._298_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._071_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._299_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._072_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._300_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._073_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._301_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._074_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._302_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._075_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._303_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._076_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._304_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._077_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._305_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._078_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._306_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._307_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._308_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._081_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._309_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._082_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._310_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._083_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._311_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._084_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._312_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._085_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._313_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._086_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._314_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._087_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._315_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._088_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._316_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._089_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._317_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._318_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._091_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._319_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._320_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._321_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._322_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._323_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._324_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._097_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._325_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._098_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._326_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._099_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._327_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._100_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._328_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._101_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._329_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._102_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._330_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._331_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._104_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._332_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._105_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._333_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._106_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._334_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._107_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._335_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._108_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._336_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._109_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._337_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._110_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._338_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._339_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._112_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._340_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._113_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._341_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._114_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._342_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._115_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._343_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._116_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._344_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._117_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._345_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._118_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._346_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._119_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._347_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._120_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._348_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._121_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._349_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._122_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._350_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._123_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._351_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._124_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._352_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._125_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._353_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._126_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._354_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._127_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._355_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._128_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._356_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._129_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._357_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._130_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._358_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._131_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._359_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._132_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._360_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._133_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._361_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._134_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._362_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._135_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._363_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._136_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._364_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._137_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._365_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._138_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._366_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._139_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._367_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._140_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._368_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._141_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._369_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._142_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._370_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._143_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._371_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._144_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._372_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._145_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._373_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._146_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._374_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._147_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._375_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._148_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._376_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._149_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._377_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._150_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._378_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._151_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._379_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._152_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._380_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._153_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._381_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._154_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._382_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._155_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._383_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._156_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._384_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._157_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._385_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._158_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._386_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._159_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._387_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._160_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._388_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._161_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._389_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._162_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._390_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._163_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._391_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._164_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._392_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._165_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._393_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._166_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._394_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._167_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._395_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._168_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._396_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._169_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._397_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._170_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._398_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._171_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._399_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._172_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._400_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._173_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._401_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._174_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._402_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._175_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._403_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._176_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._404_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._177_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._405_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._178_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._406_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._179_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._407_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._180_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._408_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._181_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._409_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._182_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._410_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._183_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._411_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._184_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._412_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._185_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._413_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._186_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._414_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._187_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._415_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._188_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._416_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._189_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._417_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._190_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._418_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._191_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._419_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._192_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._420_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._193_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._421_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._194_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._422_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._195_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._423_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._196_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._424_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._197_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._425_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._198_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._426_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._199_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._427_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._200_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._428_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._201_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._429_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._202_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._430_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._203_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._431_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._204_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._432_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._205_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._433_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._206_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._434_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._207_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._435_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._208_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._436_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._209_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._437_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._210_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._438_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._211_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._439_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._212_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._440_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._213_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._441_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._214_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._442_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._215_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._443_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._216_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._444_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._217_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._445_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._218_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._446_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._219_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._447_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._220_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._448_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._221_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._449_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._222_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._450_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem._223_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._451_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.io_oeb ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._452_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.io_out ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._453_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[0] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._454_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[1] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._455_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[2] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._456_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[3] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._457_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[4] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._458_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[5] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._459_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[6] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._460_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[7] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._461_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[8] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._462_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[9] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._463_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[10] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._464_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[11] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._465_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[12] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._466_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[13] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._467_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[14] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._468_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[15] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._469_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[16] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._470_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[17] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._471_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[18] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._472_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[19] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._473_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[20] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._474_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[21] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._475_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[22] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._476_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[23] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._477_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[24] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._478_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[25] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._479_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[26] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._480_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[27] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._481_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[28] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._482_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[29] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._483_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[30] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._484_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[31] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._485_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[32] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._486_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[33] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._487_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[34] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._488_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[35] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._489_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[36] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._490_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[37] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._491_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[38] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._492_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[39] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._493_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[40] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._494_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[41] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._495_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[42] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._496_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[43] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._497_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[44] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._498_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[45] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._499_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[46] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._500_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[47] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._501_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[48] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._502_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[49] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._503_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[50] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._504_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[51] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._505_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[52] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._506_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[53] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._507_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[54] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._508_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[55] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._509_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[56] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._510_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[57] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._511_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[58] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._512_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[59] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._513_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[60] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._514_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[61] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._515_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[62] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._516_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[63] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._517_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[64] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._518_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[65] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._519_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[66] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._520_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[67] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._521_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[68] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._522_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[69] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._523_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[70] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._524_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[71] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._525_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[72] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._526_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[73] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._527_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[74] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._528_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[75] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._529_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[76] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._530_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[77] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._531_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[78] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._532_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[79] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._533_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[80] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._534_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[81] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._535_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[82] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._536_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[83] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._537_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[84] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._538_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[85] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._539_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[86] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._540_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[87] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._541_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[88] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._542_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[89] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._543_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[90] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._544_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[91] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._545_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[92] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._546_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[93] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._547_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[94] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._548_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[95] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._549_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[96] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._550_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[97] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._551_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[98] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._552_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[99] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._553_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[100] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._554_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[101] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._555_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[102] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._556_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[103] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._557_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[104] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._558_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[105] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._559_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[106] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._560_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[107] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._561_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[108] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._562_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[109] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._563_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[110] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._564_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[111] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._565_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[112] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._566_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[113] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._567_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[114] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._568_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[115] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._569_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[116] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._570_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[117] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._571_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[118] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._572_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[119] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._573_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[120] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._574_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[121] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._575_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[122] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._576_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[123] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._577_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[124] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._578_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[125] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._579_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[126] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._580_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.la_data_out[127] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._709_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.o_irq[1] ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem._710_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.o_irq[2] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i._0609_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0000_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i._0610_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A2(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i._0001_ ));
 sky130_fd_sc_hd__nand3b_2 \efabless_subsystem.compute_controller_i._0611_  (.A_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i._0002_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i._0612_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A2(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B1_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0003_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i._0613_  (.A(\efabless_subsystem.compute_controller_i._0000_ ),
    .B(\efabless_subsystem.compute_controller_i._0001_ ),
    .C(\efabless_subsystem.compute_controller_i._0002_ ),
    .D(\efabless_subsystem.compute_controller_i._0003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0004_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0614_  (.A(\efabless_subsystem.compute_controller_i._0004_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.ctl ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i._0615_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i._0616_  (.A_N(\efabless_subsystem.compute_controller_i.acc_done_q ),
    .B(\efabless_subsystem.compute_controller_i.acc_done_q_reg.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0005_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0617_  (.A(\efabless_subsystem.compute_controller_i._0005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_done_edge ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.compute_controller_i._0618_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i._0006_ ));
 sky130_fd_sc_hd__or4bb_2 \efabless_subsystem.compute_controller_i._0619_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .C_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0007_ ));
 sky130_fd_sc_hd__or4bb_2 \efabless_subsystem.compute_controller_i._0620_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .C_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .D_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0008_ ));
 sky130_fd_sc_hd__nand3b_2 \efabless_subsystem.compute_controller_i._0621_  (.A_N(\efabless_subsystem.compute_controller_i._0006_ ),
    .B(\efabless_subsystem.compute_controller_i._0007_ ),
    .C(\efabless_subsystem.compute_controller_i._0008_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i._0622_  (.A(\efabless_subsystem.compute_controller_i._0007_ ),
    .B(\efabless_subsystem.compute_controller_i._0008_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i._0623_  (.A(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .B(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i._0009_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i._0624_  (.A1(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .A2(\efabless_subsystem.compute_controller_i._0009_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i._0625_  (.A(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i._0010_ ));
 sky130_fd_sc_hd__o211a_2 \efabless_subsystem.compute_controller_i._0626_  (.A1(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .A2(\efabless_subsystem.compute_controller_i._0009_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30.Z ),
    .C1(\efabless_subsystem.compute_controller_i._0010_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.ctl ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i._0627_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ),
    .B(\efabless_subsystem.compute_controller_i._0006_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0011_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0628_  (.A(\efabless_subsystem.compute_controller_i._0011_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i._0629_  (.A_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0012_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0630_  (.A(\efabless_subsystem.compute_controller_i._0012_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.ctl ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i._0631_  (.A_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_d[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_d[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0013_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0632_  (.A(\efabless_subsystem.compute_controller_i._0013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.o_red_params_pop ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i._0633_  (.A(\efabless_subsystem.compute_controller_i.i_acc_almost_done ),
    .B(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .C(\efabless_subsystem.compute_controller_i._0009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0014_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0634_  (.A(\efabless_subsystem.compute_controller_i._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.ctl ));
 sky130_fd_sc_hd__and4bb_2 \efabless_subsystem.compute_controller_i._0635_  (.A_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .B_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0015_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i._0636_  (.A(\efabless_subsystem.compute_controller_i.gte_709_36.Z ),
    .B(\efabless_subsystem.compute_controller_i._0015_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0016_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0637_  (.A(\efabless_subsystem.compute_controller_i._0016_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.ctl ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i._0638_  (.A(\efabless_subsystem.compute_controller_i.gte_709_36.Z ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.Z ),
    .C(\efabless_subsystem.compute_controller_i._0015_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0017_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0639_  (.A(\efabless_subsystem.compute_controller_i._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.ctl ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i._0640_  (.A(\efabless_subsystem.compute_controller_i.gte_735_31.Z ),
    .B(\efabless_subsystem.compute_controller_i.gte_734_31.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0018_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0641_  (.A(\efabless_subsystem.compute_controller_i._0018_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.ctl ));
 sky130_fd_sc_hd__o32a_2 \efabless_subsystem.compute_controller_i._0642_  (.A1(\efabless_subsystem.compute_controller_i.i_acc_almost_done ),
    .A2(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .A3(\efabless_subsystem.compute_controller_i._0009_ ),
    .B1(\efabless_subsystem.compute_controller_i._0015_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_709_36.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.ctl ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.compute_controller_i._0643_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .D_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0019_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i._0644_  (.A(\efabless_subsystem.compute_controller_i._0019_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.ctl ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.compute_controller_i._0645_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .C_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ));
 sky130_fd_sc_hd__and4bb_2 \efabless_subsystem.compute_controller_i._0646_  (.A_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i._0020_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i._0647_  (.A(\efabless_subsystem.compute_controller_i._0020_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i._0648_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1].d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i._0021_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i._0649_  (.A1(\efabless_subsystem.compute_controller_i._0021_ ),
    .A2(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2].d ),
    .B1(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.ctl ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0650_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0022_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0651_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0023_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0652_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0024_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0653_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0025_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0654_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0026_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0655_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0027_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0656_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0028_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0657_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0029_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0658_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0030_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0659_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0031_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0660_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0032_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0661_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0033_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0662_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0034_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0663_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0035_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0664_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0036_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0665_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0037_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0666_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0038_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0667_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0039_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0668_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0040_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0669_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0041_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0670_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0042_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0671_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0043_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0672_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0673_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0045_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0674_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0675_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0676_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0677_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0049_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0678_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0050_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0679_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0051_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0680_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0052_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0681_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0053_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0682_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0054_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0683_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0055_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0684_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0056_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0685_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0057_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0686_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0058_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0687_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0059_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0688_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0060_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0689_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0061_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0690_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0062_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0691_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0063_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0692_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0064_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0693_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0065_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0694_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0066_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0695_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0067_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0696_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0068_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0697_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0069_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0698_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0070_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0699_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0071_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0700_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0072_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0701_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0073_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0702_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0074_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0703_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0075_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0704_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0076_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0705_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0077_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0706_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0078_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0707_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0708_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0709_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0081_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0710_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0082_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0711_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0083_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0712_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0084_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0713_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0085_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0714_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0086_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0715_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0087_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0716_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0088_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0717_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0089_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0718_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0719_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0091_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0720_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0721_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0722_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0723_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0724_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0725_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0097_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0726_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0098_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0727_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0099_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0728_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0100_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0729_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0101_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0730_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0102_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0731_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0732_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0104_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0733_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0105_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0734_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0106_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0736_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0108_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0738_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0110_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0739_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0741_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0113_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0742_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0114_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0744_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0116_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0746_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0118_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0748_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0120_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0751_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0123_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0752_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0124_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0754_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0126_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0756_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0128_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0757_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0129_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0758_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0130_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0759_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0131_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0760_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0132_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0761_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0133_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0762_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0134_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0763_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0135_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0764_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0136_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0765_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0137_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0766_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0138_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0767_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0139_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0768_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0140_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0769_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0141_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0770_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0142_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0771_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0143_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0772_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0144_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0773_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0145_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0774_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0146_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0775_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0147_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0776_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0148_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0777_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0149_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0778_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0150_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0779_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0151_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0780_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0152_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0781_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0153_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0782_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0154_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0783_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0155_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0784_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0156_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0785_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0157_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0786_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0158_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0787_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0159_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0788_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0160_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0789_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0161_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0790_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0162_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0791_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0163_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0792_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0164_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0793_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0165_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0794_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0166_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0795_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0167_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0796_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0168_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0797_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0169_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0798_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0170_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0799_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0171_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0800_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0172_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0801_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0173_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0802_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0174_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0803_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0175_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0804_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0176_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0805_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0177_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0806_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_controller_i._0178_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0807_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0179_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0808_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0180_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0809_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0181_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0810_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0182_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0811_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0183_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0812_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0184_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0813_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0185_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0814_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0186_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0815_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0187_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0816_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0188_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0817_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0189_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0818_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0190_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0819_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0191_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0820_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0192_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0821_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0193_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0822_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0194_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0823_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0195_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0824_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0196_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0825_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0197_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0826_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0198_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0827_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0199_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0828_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0200_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0829_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0201_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0830_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0202_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0831_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0203_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0832_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0204_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0833_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0205_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0834_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0206_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0835_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0207_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0836_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0208_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0837_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0209_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0838_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0210_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0839_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0211_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0840_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0212_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0841_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0213_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0842_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0214_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0843_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0215_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0844_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0216_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0845_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0217_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0846_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0218_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0847_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0219_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0848_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0220_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0849_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0221_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0850_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0222_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0851_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0223_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0852_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0224_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0853_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0225_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0854_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0226_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0855_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0227_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0856_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0228_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0857_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0229_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0858_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0230_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0859_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0231_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0860_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0232_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0861_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0233_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0862_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0234_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0863_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0235_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0864_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0236_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0865_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0237_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0866_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0238_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0867_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0239_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0868_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0240_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0869_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0241_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0870_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0242_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0871_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0243_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0872_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0244_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0873_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0245_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0874_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0246_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0875_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0247_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0876_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0248_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0877_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0249_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0878_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0250_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0879_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0251_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0880_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0252_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0881_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0253_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0882_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0254_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0883_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0255_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0884_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0256_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0885_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0257_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0886_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0258_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0887_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0259_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0888_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0260_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0889_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0261_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0890_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0262_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0891_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0263_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0892_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0264_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0893_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0265_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0894_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0266_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0895_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0267_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0896_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0268_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0897_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0269_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0898_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0270_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0899_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0271_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0900_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0272_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0901_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0273_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0902_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0274_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0903_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0275_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0904_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0276_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0905_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0277_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0906_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0278_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0907_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0279_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0908_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0280_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0909_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0281_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0910_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0282_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0911_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0283_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0912_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0284_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0913_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0285_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0914_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0286_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0915_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0287_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0916_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0288_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0917_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0289_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0918_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0290_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0919_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0291_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0920_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0292_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0921_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0293_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0922_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0294_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0923_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0295_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0924_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0296_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0925_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0297_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0926_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0298_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0927_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0299_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0928_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0300_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0929_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0301_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0930_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0302_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0931_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0303_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0932_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0304_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0933_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0305_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0934_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0306_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0935_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0307_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0936_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0308_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0937_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0309_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0938_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0310_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0939_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0311_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0940_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0312_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0941_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0313_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0942_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0314_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0943_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0315_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0944_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0316_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0945_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0317_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0946_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0318_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0947_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0319_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0948_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0320_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0949_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0321_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0950_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0322_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0951_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0323_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0952_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0324_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0953_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0325_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0954_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0326_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0955_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0327_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0956_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0328_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0957_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0329_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0958_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0330_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0959_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0331_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0960_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0332_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0961_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0333_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0962_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0334_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0963_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0335_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0964_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0336_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0965_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0337_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0966_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0338_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0967_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0339_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0968_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0340_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0969_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0341_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0970_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0342_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0971_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0343_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0972_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0344_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0973_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0345_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0974_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0346_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0975_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0347_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0976_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0348_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0977_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0349_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0978_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0350_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0979_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0351_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0980_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0352_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0981_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0353_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0982_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0354_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0983_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0355_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0984_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0356_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0985_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0357_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0986_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0358_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0987_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0359_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0988_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0360_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0989_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0361_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0990_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0362_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0991_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0363_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0992_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0364_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0993_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0365_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0994_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0366_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0995_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0367_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0996_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0368_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0997_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0369_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._0999_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0371_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1000_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0372_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1001_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0373_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1002_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0374_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1003_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0375_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1004_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0376_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1005_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0377_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1006_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0378_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1007_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0379_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1008_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0380_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1009_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0381_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1010_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0382_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1011_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0383_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1012_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0384_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1013_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0385_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1014_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0386_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1015_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0387_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1016_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0388_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1017_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0389_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1018_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0390_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1019_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0391_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1020_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0392_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1021_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0393_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1022_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0394_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1023_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0395_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1024_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0396_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1025_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0397_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1029_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0401_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1030_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0402_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1031_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0403_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1035_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0407_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1036_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0408_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1040_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0412_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1041_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0413_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1042_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0414_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1046_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0418_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1047_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0419_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1048_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0420_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1051_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0423_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1052_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0424_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1055_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0427_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1058_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0430_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1059_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0431_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1063_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0435_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1064_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0436_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1067_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0439_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1068_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0440_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1071_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0443_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1072_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0444_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1075_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0447_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1076_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0448_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1078_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0450_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1080_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0452_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1083_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0455_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1085_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0457_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1086_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0458_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1088_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0460_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1089_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0461_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1090_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0462_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1091_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0463_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1092_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0464_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1093_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0465_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1094_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0466_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1095_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0467_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1096_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0468_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1097_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0469_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1098_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0470_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1099_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0471_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1100_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0472_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1101_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0473_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1102_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0474_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1103_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0475_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1104_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0476_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1105_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0477_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1106_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0478_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1107_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0479_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1108_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0480_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1109_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0481_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1110_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0482_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1111_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0483_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1112_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0484_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1113_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0485_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1114_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0486_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1115_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0487_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1116_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0488_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1117_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0489_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1118_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0490_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1119_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0491_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1120_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0492_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1121_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0493_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1122_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0494_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1123_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0495_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1124_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0496_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1125_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0497_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1126_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0498_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1127_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0499_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1128_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0500_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1129_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0501_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1130_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0502_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1131_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0503_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1132_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0504_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1133_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0505_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1134_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0506_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1135_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0507_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1136_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0508_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1137_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0509_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1138_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0510_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1139_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0511_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1140_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0512_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1141_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0513_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1142_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0514_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1143_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0515_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1144_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0516_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1145_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0517_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1146_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0518_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1147_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0519_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1148_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0520_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1149_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0521_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1150_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0522_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1151_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0523_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1152_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0524_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1153_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0525_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1154_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0526_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1155_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0527_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1156_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0528_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1157_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0529_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1158_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0530_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1159_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0531_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1160_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0532_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1161_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0533_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1162_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0534_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1163_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0535_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1164_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0536_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1165_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0537_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1166_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0538_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1167_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0539_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1168_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0540_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1169_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0541_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1170_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0542_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1171_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0543_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1172_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0544_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1173_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0545_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1174_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0546_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1175_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0547_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1176_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0548_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1177_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0549_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1178_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0550_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1179_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0551_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1180_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0552_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1181_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0553_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1182_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0554_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1183_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0555_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1184_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0556_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1185_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0557_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1186_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0558_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1187_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0559_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1188_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0560_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1189_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0561_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1190_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0562_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1191_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0563_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1192_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0564_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1193_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0565_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1194_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0566_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1195_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0567_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1196_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0568_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1197_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0569_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1198_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0570_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1199_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0571_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1200_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0572_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1201_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0573_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1202_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0574_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1203_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0575_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1204_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0576_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1205_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0577_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1206_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0578_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1207_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0579_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1208_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0580_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1209_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0581_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1210_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0582_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1211_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0583_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1212_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0584_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1213_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0585_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1214_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0586_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1215_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0587_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1216_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0588_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1217_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0589_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1218_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0590_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1219_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0591_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1220_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0592_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1221_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0593_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1222_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0594_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1223_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0595_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1224_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0596_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1225_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0597_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1226_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0598_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1227_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0599_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1228_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0600_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1229_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0601_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1230_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0602_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1231_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0603_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1232_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0604_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1233_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0605_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1234_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0606_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1235_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0607_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_controller_i._1236_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_controller_i._0608_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0179_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[0] ),
    .S(\efabless_subsystem.compute_controller_i._0022_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0180_ ),
    .S(\efabless_subsystem.compute_controller_i._0181_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0182_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[10] ),
    .S(\efabless_subsystem.compute_controller_i._0023_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0183_ ),
    .S(\efabless_subsystem.compute_controller_i._0184_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0185_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[11] ),
    .S(\efabless_subsystem.compute_controller_i._0024_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0186_ ),
    .S(\efabless_subsystem.compute_controller_i._0187_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0188_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[12] ),
    .S(\efabless_subsystem.compute_controller_i._0025_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0189_ ),
    .S(\efabless_subsystem.compute_controller_i._0190_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0191_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[13] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[13] ),
    .S(\efabless_subsystem.compute_controller_i._0026_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0192_ ),
    .S(\efabless_subsystem.compute_controller_i._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[13] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[13]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0194_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[14] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[14] ),
    .S(\efabless_subsystem.compute_controller_i._0027_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0195_ ),
    .S(\efabless_subsystem.compute_controller_i._0196_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[14] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[14]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0197_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[15] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[15] ),
    .S(\efabless_subsystem.compute_controller_i._0028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0198_ ),
    .S(\efabless_subsystem.compute_controller_i._0199_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[15] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[15]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0200_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[1] ),
    .S(\efabless_subsystem.compute_controller_i._0029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0201_ ),
    .S(\efabless_subsystem.compute_controller_i._0202_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0203_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[2] ),
    .S(\efabless_subsystem.compute_controller_i._0030_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0204_ ),
    .S(\efabless_subsystem.compute_controller_i._0205_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0206_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[3] ),
    .S(\efabless_subsystem.compute_controller_i._0031_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0207_ ),
    .S(\efabless_subsystem.compute_controller_i._0208_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0209_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[4] ),
    .S(\efabless_subsystem.compute_controller_i._0032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0210_ ),
    .S(\efabless_subsystem.compute_controller_i._0211_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0212_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[5] ),
    .S(\efabless_subsystem.compute_controller_i._0033_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0213_ ),
    .S(\efabless_subsystem.compute_controller_i._0214_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0215_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[6] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[6] ),
    .S(\efabless_subsystem.compute_controller_i._0034_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0216_ ),
    .S(\efabless_subsystem.compute_controller_i._0217_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[6] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[7] ),
    .S(\efabless_subsystem.compute_controller_i._0035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0219_ ),
    .S(\efabless_subsystem.compute_controller_i._0220_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[8] ),
    .S(\efabless_subsystem.compute_controller_i._0036_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0222_ ),
    .S(\efabless_subsystem.compute_controller_i._0223_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0224_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[9] ),
    .S(\efabless_subsystem.compute_controller_i._0037_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0225_ ),
    .S(\efabless_subsystem.compute_controller_i._0226_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_done_q_reg._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_done_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_done_q_reg._08_  (.A(\efabless_subsystem.compute_controller_i.acc_done_q_reg._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0227_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_done_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_done_q_reg._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_done_q ),
    .A1(\efabless_subsystem.compute_controller_i.acc_done_q_reg.d ),
    .S(\efabless_subsystem.compute_controller_i._0038_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_done_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_done_q_reg._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_done_q_reg._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0228_ ),
    .S(\efabless_subsystem.compute_controller_i._0229_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_done_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_done_q_reg._11_  (.A(\efabless_subsystem.compute_controller_i.acc_done_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_done_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_done_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_done_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_done_q_reg._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_done_q_reg._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_done_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_done_q_reg._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_done_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_done_q ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_done_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0230_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q ),
    .A1(\efabless_subsystem.compute_controller_i.acc_pos_cnt_d ),
    .S(\efabless_subsystem.compute_controller_i._0039_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0231_ ),
    .S(\efabless_subsystem.compute_controller_i._0232_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q ),
    .Q_N(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_143_38._0_  (.A(\efabless_subsystem.compute_controller_i._0040_ ),
    .B(\efabless_subsystem.compute_controller_i.add_143_38.A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_143_38.Z ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_157_42._0_  (.A(\efabless_subsystem.compute_controller_i._0041_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_157_42.Z ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_163_38._3_  (.A(\efabless_subsystem.compute_controller_i._0042_ ),
    .B(\efabless_subsystem.compute_controller_i.add_163_38.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_163_38._0_ ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_163_38._4_  (.A(\efabless_subsystem.compute_controller_i.add_163_38.A[1] ),
    .B(\efabless_subsystem.compute_controller_i.add_163_38._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_163_38.Z[1] ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.add_163_38._5_  (.A(\efabless_subsystem.compute_controller_i._0042_ ),
    .B(\efabless_subsystem.compute_controller_i.add_163_38.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_163_38._1_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_163_38._6_  (.A(\efabless_subsystem.compute_controller_i.add_163_38._0_ ),
    .B(\efabless_subsystem.compute_controller_i.add_163_38._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_163_38._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_163_38._7_  (.A(\efabless_subsystem.compute_controller_i.add_163_38._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_163_38.Z[0] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_175_34._24_  (.A(\efabless_subsystem.compute_controller_i._0043_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._00_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.add_175_34._25_  (.A1(\efabless_subsystem.compute_controller_i._0043_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .B1(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34._01_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_175_34._26_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._00_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34.Z[1] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_175_34._27_  (.A(\efabless_subsystem.compute_controller_i._0043_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .D(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_175_34._28_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_175_34._29_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._02_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34.Z[2] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_175_34._30_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34._04_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_175_34._31_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_175_34._32_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._04_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34.Z[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_175_34._33_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[4] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_175_34._34_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._06_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_175_34._35_  (.A1(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .A3(\efabless_subsystem.compute_controller_i.add_175_34._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._07_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.add_175_34._36_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34._06_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_175_34._37_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_175_34._38_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[6] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_175_34._39_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_175_34._40_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34._02_ ),
    .D(\efabless_subsystem.compute_controller_i.add_175_34._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_175_34._41_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._11_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_175_34._42_  (.A1(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34._02_ ),
    .A3(\efabless_subsystem.compute_controller_i.add_175_34._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._12_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.add_175_34._43_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_175_34._44_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_175_34._45_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[8] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_175_34._46_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._14_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.add_175_34._47_  (.A1(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34._15_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_175_34._48_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._14_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34.Z[9] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_175_34._49_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .D(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._16_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.compute_controller_i.add_175_34._50_  (.A1(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.add_175_34._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[10] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_175_34._51_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .D(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._17_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_175_34._52_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34._18_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.add_175_34._53_  (.A1(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_175_34._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[11] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_175_34._54_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34.Z[12] ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_175_34._55_  (.A1(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .A2(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .A3(\efabless_subsystem.compute_controller_i.add_175_34._17_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._19_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_175_34._56_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._20_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_175_34._57_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34._21_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_175_34._58_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._19_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._22_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_175_34._59_  (.A(\efabless_subsystem.compute_controller_i.add_175_34._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[13] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_175_34._60_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_175_34.Z[14] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_175_34._61_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._11_ ),
    .C(\efabless_subsystem.compute_controller_i.add_175_34._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34._23_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_175_34._62_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34._23_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[15] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_175_34._63_  (.A(\efabless_subsystem.compute_controller_i._0043_ ),
    .B(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_175_34.Z[0] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_185_30._24_  (.A(\efabless_subsystem.compute_controller_i._0044_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .C(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._00_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.add_185_30._25_  (.A1(\efabless_subsystem.compute_controller_i._0044_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30._01_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_185_30._26_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._00_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30.Z[1] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_185_30._27_  (.A(\efabless_subsystem.compute_controller_i._0044_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .C(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_185_30._28_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_185_30._29_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._02_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30.Z[2] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_185_30._30_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30._04_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_185_30._31_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_185_30._32_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._04_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30.Z[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_185_30._33_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[4] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_185_30._34_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.add_185_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._06_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_185_30._35_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .A3(\efabless_subsystem.compute_controller_i.add_185_30._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._07_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.add_185_30._36_  (.A_N(\efabless_subsystem.compute_controller_i.add_185_30._06_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_185_30._37_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_185_30._38_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[6] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[6] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_185_30._39_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.acc_cnt_q[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_185_30._40_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .C(\efabless_subsystem.compute_controller_i.add_185_30._02_ ),
    .D(\efabless_subsystem.compute_controller_i.add_185_30._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_185_30._41_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._11_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_185_30._42_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.add_185_30._02_ ),
    .A3(\efabless_subsystem.compute_controller_i.add_185_30._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._12_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.add_185_30._43_  (.A_N(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_185_30._44_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_185_30._45_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[8] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_185_30._46_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._14_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.add_185_30._47_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .A2(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30._15_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_185_30._48_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._14_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30.Z[9] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_185_30._49_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .D(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._16_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.compute_controller_i.add_185_30._50_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .A2(\efabless_subsystem.compute_controller_i.add_185_30._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.add_185_30._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[10] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_185_30._51_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .D(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._17_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_185_30._52_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30._18_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.add_185_30._53_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .A2(\efabless_subsystem.compute_controller_i.add_185_30._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_185_30._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[11] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_185_30._54_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30.Z[12] ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_185_30._55_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .A2(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .A3(\efabless_subsystem.compute_controller_i.add_185_30._17_ ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_q[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._19_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_185_30._56_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[13] ),
    .C(\efabless_subsystem.compute_controller_i.add_185_30._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._20_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_185_30._57_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30._21_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_185_30._58_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._19_ ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._22_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_185_30._59_  (.A(\efabless_subsystem.compute_controller_i.add_185_30._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[13] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_185_30._60_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[14] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_185_30.Z[14] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_185_30._61_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[14] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._11_ ),
    .C(\efabless_subsystem.compute_controller_i.add_185_30._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30._23_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_185_30._62_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[15] ),
    .B(\efabless_subsystem.compute_controller_i.add_185_30._23_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[15] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_185_30._63_  (.A(\efabless_subsystem.compute_controller_i._0044_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_185_30.Z[0] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_200_30._24_  (.A(\efabless_subsystem.compute_controller_i._0045_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._00_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.add_200_30._25_  (.A1(\efabless_subsystem.compute_controller_i._0045_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30._01_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_200_30._26_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._00_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30.Z[1] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_200_30._27_  (.A(\efabless_subsystem.compute_controller_i._0045_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .D(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_200_30._28_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_200_30._29_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._02_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30.Z[2] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_200_30._30_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30._04_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_200_30._31_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_200_30._32_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._04_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30.Z[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_200_30._33_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[4] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_200_30._34_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._06_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_200_30._35_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .A3(\efabless_subsystem.compute_controller_i.add_200_30._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._07_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.add_200_30._36_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30._06_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_200_30._37_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_200_30._38_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[6] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_200_30._39_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_200_30._40_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30._02_ ),
    .D(\efabless_subsystem.compute_controller_i.add_200_30._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_200_30._41_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._11_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_200_30._42_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30._02_ ),
    .A3(\efabless_subsystem.compute_controller_i.add_200_30._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._12_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.add_200_30._43_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_200_30._44_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_200_30._45_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[8] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_200_30._46_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._14_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.add_200_30._47_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30._15_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.add_200_30._48_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._14_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30.Z[9] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_200_30._49_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .D(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._16_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.compute_controller_i.add_200_30._50_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.add_200_30._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[10] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.compute_controller_i.add_200_30._51_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .D(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._17_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_200_30._52_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30._18_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.add_200_30._53_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[11] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_200_30._54_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30.Z[12] ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.add_200_30._55_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .A3(\efabless_subsystem.compute_controller_i.add_200_30._17_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._19_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_200_30._56_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._20_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.add_200_30._57_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30._21_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.add_200_30._58_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._19_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._22_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.add_200_30._59_  (.A(\efabless_subsystem.compute_controller_i.add_200_30._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[13] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.add_200_30._60_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.add_200_30.Z[14] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.add_200_30._61_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._11_ ),
    .C(\efabless_subsystem.compute_controller_i.add_200_30._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30._23_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_200_30._62_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30._23_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[15] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.add_200_30._63_  (.A(\efabless_subsystem.compute_controller_i._0045_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.add_200_30.Z[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0233_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].d ),
    .S(\efabless_subsystem.compute_controller_i._0046_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0234_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0235_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1].d ),
    .S(\efabless_subsystem.compute_controller_i._0047_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0236_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0237_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2].d ),
    .S(\efabless_subsystem.compute_controller_i._0048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0238_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0239_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0].d ),
    .S(\efabless_subsystem.compute_controller_i._0049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0240_ ),
    .S(\efabless_subsystem.compute_controller_i._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0242_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10].d ),
    .S(\efabless_subsystem.compute_controller_i._0050_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0243_ ),
    .S(\efabless_subsystem.compute_controller_i._0244_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0245_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11].d ),
    .S(\efabless_subsystem.compute_controller_i._0051_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0246_ ),
    .S(\efabless_subsystem.compute_controller_i._0247_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0248_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12].d ),
    .S(\efabless_subsystem.compute_controller_i._0052_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0249_ ),
    .S(\efabless_subsystem.compute_controller_i._0250_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13].d ),
    .S(\efabless_subsystem.compute_controller_i._0053_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0252_ ),
    .S(\efabless_subsystem.compute_controller_i._0253_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0254_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14].d ),
    .S(\efabless_subsystem.compute_controller_i._0054_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0255_ ),
    .S(\efabless_subsystem.compute_controller_i._0256_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0257_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15].d ),
    .S(\efabless_subsystem.compute_controller_i._0055_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0258_ ),
    .S(\efabless_subsystem.compute_controller_i._0259_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0260_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1].d ),
    .S(\efabless_subsystem.compute_controller_i._0056_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0261_ ),
    .S(\efabless_subsystem.compute_controller_i._0262_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0263_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2].d ),
    .S(\efabless_subsystem.compute_controller_i._0057_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0264_ ),
    .S(\efabless_subsystem.compute_controller_i._0265_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0266_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3].d ),
    .S(\efabless_subsystem.compute_controller_i._0058_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0267_ ),
    .S(\efabless_subsystem.compute_controller_i._0268_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0269_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4].d ),
    .S(\efabless_subsystem.compute_controller_i._0059_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0270_ ),
    .S(\efabless_subsystem.compute_controller_i._0271_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0272_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5].d ),
    .S(\efabless_subsystem.compute_controller_i._0060_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0273_ ),
    .S(\efabless_subsystem.compute_controller_i._0274_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0275_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6].d ),
    .S(\efabless_subsystem.compute_controller_i._0061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0276_ ),
    .S(\efabless_subsystem.compute_controller_i._0277_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0278_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7].d ),
    .S(\efabless_subsystem.compute_controller_i._0062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0279_ ),
    .S(\efabless_subsystem.compute_controller_i._0280_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0281_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8].d ),
    .S(\efabless_subsystem.compute_controller_i._0063_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0282_ ),
    .S(\efabless_subsystem.compute_controller_i._0283_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._08_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0284_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._09_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9].d ),
    .S(\efabless_subsystem.compute_controller_i._0064_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._10_  (.A0(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0285_ ),
    .S(\efabless_subsystem.compute_controller_i._0286_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._11_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .Q_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0287_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_163_38.A[0] ),
    .A1(\efabless_subsystem.compute_controller_i.aux_pos_cnt_d[0] ),
    .S(\efabless_subsystem.compute_controller_i._0065_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0288_ ),
    .S(\efabless_subsystem.compute_controller_i._0289_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_163_38.A[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0290_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_163_38.A[1] ),
    .A1(\efabless_subsystem.compute_controller_i.aux_pos_cnt_d[1] ),
    .S(\efabless_subsystem.compute_controller_i._0066_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0291_ ),
    .S(\efabless_subsystem.compute_controller_i._0292_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_163_38.A[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.aux_pos_cnt_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0293_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].d ),
    .S(\efabless_subsystem.compute_controller_i._0067_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0294_ ),
    .S(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0295_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1].d ),
    .S(\efabless_subsystem.compute_controller_i._0068_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0296_ ),
    .S(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._08_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0297_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._09_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2].d ),
    .S(\efabless_subsystem.compute_controller_i._0069_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._10_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0298_ ),
    .S(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._11_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .Q_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._08_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0299_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._09_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3].d ),
    .S(\efabless_subsystem.compute_controller_i._0070_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._10_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0300_ ),
    .S(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._11_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .Q_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3]._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._14_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._15_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.ctl_375_11._16_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._02_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.compute_controller_i.ctl_375_11._17_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .B(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[11] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.ctl_375_11._18_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_375_11._03_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.compute_controller_i.ctl_375_11._19_  (.A_N(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .B(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._04_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._20_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[10] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.compute_controller_i.ctl_375_11._21_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .D_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._05_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctl_375_11._22_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[9] ));
 sky130_fd_sc_hd__and4bb_2 \efabless_subsystem.compute_controller_i.ctl_375_11._23_  (.A_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B_N(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._24_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[8] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.compute_controller_i.ctl_375_11._25_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .D_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._07_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctl_375_11._26_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[7] ));
 sky130_fd_sc_hd__and4bb_2 \efabless_subsystem.compute_controller_i.ctl_375_11._27_  (.A_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .B_N(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._28_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[6] ));
 sky130_fd_sc_hd__and4bb_2 \efabless_subsystem.compute_controller_i.ctl_375_11._29_  (.A_N(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .B_N(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._09_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._30_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[5] ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.compute_controller_i.ctl_375_11._31_  (.A_N(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .B(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .C(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._32_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[4] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.compute_controller_i.ctl_375_11._33_  (.A_N(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .B(\efabless_subsystem.compute_controller_i.ctl_375_11._03_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._11_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._34_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[3] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.ctl_375_11._35_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .B(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._12_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._36_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[2] ));
 sky130_fd_sc_hd__and4bb_2 \efabless_subsystem.compute_controller_i.ctl_375_11._37_  (.A_N(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .B_N(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .C(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .D(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_375_11._38_  (.A(\efabless_subsystem.compute_controller_i.ctl_375_11._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[1] ));
 sky130_fd_sc_hd__o211a_2 \efabless_subsystem.compute_controller_i.ctl_375_11._39_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11._01_ ),
    .B1(\efabless_subsystem.compute_controller_i.ctl_375_11._02_ ),
    .C1(\efabless_subsystem.compute_controller_i.ctl_375_11._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[0] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.compute_controller_i.ctl_775_11._03_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .C(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[6] ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.compute_controller_i.ctl_775_11._04_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .C_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[5] ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.compute_controller_i.ctl_775_11._05_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .C_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[4] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.compute_controller_i.ctl_775_11._06_  (.A_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .C(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_775_11._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_775_11._07_  (.A(\efabless_subsystem.compute_controller_i.ctl_775_11._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[3] ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.compute_controller_i.ctl_775_11._08_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .C_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[2] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.compute_controller_i.ctl_775_11._09_  (.A_N(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .C(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_775_11._01_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_775_11._10_  (.A(\efabless_subsystem.compute_controller_i.ctl_775_11._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[1] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.ctl_775_11._11_  (.A(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_775_11._02_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_775_11._12_  (.A(\efabless_subsystem.compute_controller_i.ctl_775_11._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[0] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._3_  (.A(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .B(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[3] ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._4_  (.A_N(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .B(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._5_  (.A(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[2] ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._6_  (.A_N(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .B(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._7_  (.A(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[1] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._8_  (.A(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .B(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._1_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._9_  (.A(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0301_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[0] ),
    .S(\efabless_subsystem.compute_controller_i._0071_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0302_ ),
    .S(\efabless_subsystem.compute_controller_i._0303_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0304_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[10] ),
    .S(\efabless_subsystem.compute_controller_i._0072_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0305_ ),
    .S(\efabless_subsystem.compute_controller_i._0306_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0307_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[11] ),
    .S(\efabless_subsystem.compute_controller_i._0073_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0308_ ),
    .S(\efabless_subsystem.compute_controller_i._0309_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0310_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[12] ),
    .S(\efabless_subsystem.compute_controller_i._0074_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0311_ ),
    .S(\efabless_subsystem.compute_controller_i._0312_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0313_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[13] ),
    .S(\efabless_subsystem.compute_controller_i._0075_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0314_ ),
    .S(\efabless_subsystem.compute_controller_i._0315_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[13]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0316_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[14] ),
    .S(\efabless_subsystem.compute_controller_i._0076_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0317_ ),
    .S(\efabless_subsystem.compute_controller_i._0318_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[14]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0319_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[15] ),
    .S(\efabless_subsystem.compute_controller_i._0077_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0320_ ),
    .S(\efabless_subsystem.compute_controller_i._0321_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[15]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0322_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[1] ),
    .S(\efabless_subsystem.compute_controller_i._0078_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0323_ ),
    .S(\efabless_subsystem.compute_controller_i._0324_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0325_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[2] ),
    .S(\efabless_subsystem.compute_controller_i._0079_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0326_ ),
    .S(\efabless_subsystem.compute_controller_i._0327_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0328_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[3] ),
    .S(\efabless_subsystem.compute_controller_i._0080_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0329_ ),
    .S(\efabless_subsystem.compute_controller_i._0330_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0331_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[4] ),
    .S(\efabless_subsystem.compute_controller_i._0081_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0332_ ),
    .S(\efabless_subsystem.compute_controller_i._0333_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0334_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[5] ),
    .S(\efabless_subsystem.compute_controller_i._0082_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0335_ ),
    .S(\efabless_subsystem.compute_controller_i._0336_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0337_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[6] ),
    .S(\efabless_subsystem.compute_controller_i._0083_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0338_ ),
    .S(\efabless_subsystem.compute_controller_i._0339_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0340_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[7] ),
    .S(\efabless_subsystem.compute_controller_i._0084_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0341_ ),
    .S(\efabless_subsystem.compute_controller_i._0342_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0343_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[8] ),
    .S(\efabless_subsystem.compute_controller_i._0085_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0344_ ),
    .S(\efabless_subsystem.compute_controller_i._0345_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._08_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0346_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .A1(\efabless_subsystem.compute_controller_i.ctx_cnt_d[9] ),
    .S(\efabless_subsystem.compute_controller_i._0086_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._10_  (.A0(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0347_ ),
    .S(\efabless_subsystem.compute_controller_i._0348_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._11_  (.A(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .Q_N(\efabless_subsystem.compute_controller_i.ctx_cnt_q_reg[9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gt_269_32._07_  (.A(\efabless_subsystem.compute_controller_i._0087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gt_269_32._00_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gt_269_32._08_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .A2(\efabless_subsystem.compute_controller_i.gt_269_32._00_ ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .C1(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gt_269_32._09_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gt_269_32._10_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[1] ),
    .D(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32._03_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gt_269_32._11_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .D(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32._04_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gt_269_32._12_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32._02_ ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32._03_ ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32._05_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gt_269_32._13_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32._01_ ),
    .D(\efabless_subsystem.compute_controller_i.gt_269_32._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.gt_269_32._14_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gt_269_32.Z ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.gte_255_34._1_  (.A(\efabless_subsystem.compute_controller_i.add_143_38.A ),
    .B_N(\efabless_subsystem.compute_controller_i._0088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_255_34._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.gte_255_34._2_  (.A(\efabless_subsystem.compute_controller_i.gte_255_34._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_255_34.Z ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.gte_262_34._1_  (.A(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q ),
    .B_N(\efabless_subsystem.compute_controller_i._0089_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_262_34._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.gte_262_34._2_  (.A(\efabless_subsystem.compute_controller_i.gte_262_34._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_262_34.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._44_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._00_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._45_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._46_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._02_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_286_30._47_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_d[1] ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_d[0] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._48_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._04_ ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.gte_286_30._49_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[3] ),
    .B_N(\efabless_subsystem.compute_controller_i.gte_286_30.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._05_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.gte_286_30._50_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._04_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_d[2] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._01_ ),
    .B2(\efabless_subsystem.compute_controller_i.acc_cnt_d[1] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._06_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.gte_286_30._51_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30._04_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_d[2] ),
    .C(\efabless_subsystem.compute_controller_i.gte_286_30._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._07_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_286_30._52_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_d[3] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._00_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._03_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._08_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._53_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._09_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._54_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._55_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._11_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_286_30._56_  (.A_N(\efabless_subsystem.compute_controller_i.acc_cnt_d[7] ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._12_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_286_30._57_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._10_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._11_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._13_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_286_30._58_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._14_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._59_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._15_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_286_30._60_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._11_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._15_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._16_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._61_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._17_ ));
 sky130_fd_sc_hd__o2bb2a_2 \efabless_subsystem.compute_controller_i.gte_286_30._62_  (.A1_N(\efabless_subsystem.compute_controller_i.gte_286_30._17_ ),
    .A2_N(\efabless_subsystem.compute_controller_i.acc_cnt_d[4] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._18_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_286_30._63_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._11_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._19_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_286_30._64_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._12_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._18_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._20_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.gte_286_30._65_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._08_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.gte_286_30._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._21_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._66_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._22_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._67_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._23_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._68_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._24_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._69_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._25_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_286_30._70_  (.A_N(\efabless_subsystem.compute_controller_i.acc_cnt_d[15] ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._26_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_286_30._71_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[13] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._24_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._25_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[14] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._26_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._27_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_286_30._72_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._28_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._73_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._29_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.gte_286_30._74_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30._29_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_d[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._30_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._75_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._31_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_286_30._76_  (.A_N(\efabless_subsystem.compute_controller_i.acc_cnt_d[11] ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._32_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_286_30._77_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._31_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[10] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._33_ ));
 sky130_fd_sc_hd__o2111a_2 \efabless_subsystem.compute_controller_i.gte_286_30._78_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_d[8] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._28_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._30_ ),
    .D1(\efabless_subsystem.compute_controller_i.gte_286_30._33_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._34_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.compute_controller_i.gte_286_30._79_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30._31_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[10] ),
    .C(\efabless_subsystem.compute_controller_i.gte_286_30._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._35_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_286_30._80_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_d[8] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._29_ ),
    .B2(\efabless_subsystem.compute_controller_i.acc_cnt_d[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._36_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._81_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._37_ ));
 sky130_fd_sc_hd__a32o_2 \efabless_subsystem.compute_controller_i.gte_286_30._82_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._30_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._33_ ),
    .A3(\efabless_subsystem.compute_controller_i.gte_286_30._36_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._37_ ),
    .B2(\efabless_subsystem.compute_controller_i.acc_cnt_d[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._38_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_286_30._83_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._35_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._38_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._28_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._39_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_286_30._84_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_d[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._40_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_286_30._85_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._25_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[14] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._40_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._41_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_286_30._86_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30._42_ ));
 sky130_fd_sc_hd__o22ai_2 \efabless_subsystem.compute_controller_i.gte_286_30._87_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._26_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._41_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._42_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_286_30._43_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_286_30._88_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30._21_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30._34_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30._39_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_286_30._43_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_286_30.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._050_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._000_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._051_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._001_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_678_56._052_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[2] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._000_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._001_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._002_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._053_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._003_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._054_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._004_ ));
 sky130_fd_sc_hd__o211a_2 \efabless_subsystem.compute_controller_i.gte_678_56._055_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[1] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._003_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._004_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56.B[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._005_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_678_56._056_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[2] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._000_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[1] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56._003_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56._005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._006_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._057_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._007_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.gte_678_56._058_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[5] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._008_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._059_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._009_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._060_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._010_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_678_56._061_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._009_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[6] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._010_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._011_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._062_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._012_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_678_56._063_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._012_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._001_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._013_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_678_56._064_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56._008_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56._011_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56._013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._014_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_678_56._065_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._002_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._006_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._015_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_678_56._066_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._010_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[7] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._016_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_678_56._067_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._010_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[7] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._016_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56.B[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._017_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_678_56._068_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._012_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[5] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._018_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_678_56._069_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56._008_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56._011_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56._018_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._019_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._070_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._020_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._071_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._021_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._072_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._022_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_678_56._073_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._023_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._074_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._024_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_678_56._075_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._025_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_678_56._076_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._026_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_678_56._077_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._027_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.gte_678_56._078_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._024_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._025_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56._026_ ),
    .D1(\efabless_subsystem.compute_controller_i.gte_678_56._027_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._028_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_678_56._079_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._022_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[10] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._023_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56._028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._029_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_678_56._080_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._020_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56._021_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56._029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._030_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.gte_678_56._081_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._015_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._017_ ),
    .A3(\efabless_subsystem.compute_controller_i.gte_678_56._019_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._030_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._031_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_678_56._082_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._020_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56._021_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._032_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_678_56._083_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[9] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._021_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._033_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._084_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._034_ ));
 sky130_fd_sc_hd__or3b_2 \efabless_subsystem.compute_controller_i.gte_678_56._085_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[10] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56._023_ ),
    .C_N(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._035_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_678_56._086_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._034_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[11] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._036_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._087_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._037_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._088_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._038_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_678_56._089_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._037_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[14] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._038_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._039_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_678_56._090_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56._040_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_678_56._091_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._024_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56._040_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._041_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_678_56._092_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56._025_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56._026_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56._027_ ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56._041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._042_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.gte_678_56._093_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._028_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._036_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._039_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56._027_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56._042_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._043_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_678_56._094_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._029_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._033_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._044_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_678_56._095_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[25] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[24] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[27] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._045_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_678_56._096_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[21] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[20] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[23] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._046_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_678_56._097_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[17] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[16] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[19] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._047_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_678_56._098_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[29] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[28] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._048_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_678_56._099_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56._046_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56._047_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56._048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56._049_ ));
 sky130_fd_sc_hd__a211oi_2 \efabless_subsystem.compute_controller_i.gte_678_56._100_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56._031_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56._044_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56._045_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56._049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._050_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._000_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._051_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._001_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_688_48._052_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[2] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._000_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._001_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._002_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._053_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._003_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._054_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._004_ ));
 sky130_fd_sc_hd__o211a_2 \efabless_subsystem.compute_controller_i.gte_688_48._055_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[1] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._003_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._004_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48.B[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._005_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_688_48._056_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[2] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._000_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48.B[1] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48._003_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48._005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._006_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._057_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._007_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.gte_688_48._058_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[5] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._008_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._059_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._009_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._060_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._010_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_688_48._061_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._009_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[6] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._010_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._011_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._062_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._012_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_688_48._063_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._012_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._001_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._013_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_688_48._064_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48._008_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48._011_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48._013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._014_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_688_48._065_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._002_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._006_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._015_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_688_48._066_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._010_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[7] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._016_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_688_48._067_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._010_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[7] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._016_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48.B[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._017_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_688_48._068_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._012_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48.B[5] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._018_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_688_48._069_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48._008_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48._011_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48._018_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._019_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._070_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._020_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._071_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._021_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._072_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._022_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_688_48._073_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._023_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._074_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._024_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_688_48._075_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._025_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_688_48._076_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._026_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_688_48._077_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._027_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.gte_688_48._078_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._024_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._025_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48._026_ ),
    .D1(\efabless_subsystem.compute_controller_i.gte_688_48._027_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._028_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_688_48._079_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._022_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[10] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._023_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48._028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._029_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_688_48._080_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._020_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48._021_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48._029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._030_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.gte_688_48._081_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._015_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._017_ ),
    .A3(\efabless_subsystem.compute_controller_i.gte_688_48._019_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._030_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._031_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_688_48._082_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._020_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48._021_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._032_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_688_48._083_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48.B[9] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._021_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._033_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._084_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._034_ ));
 sky130_fd_sc_hd__or3b_2 \efabless_subsystem.compute_controller_i.gte_688_48._085_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[10] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48._023_ ),
    .C_N(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._035_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_688_48._086_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._034_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[11] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._036_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._087_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._037_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._088_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._038_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_688_48._089_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._037_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[14] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._038_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._039_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_688_48._090_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48._040_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_688_48._091_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._024_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48._040_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._041_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_688_48._092_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48._025_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48._026_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48._027_ ),
    .D(\efabless_subsystem.compute_controller_i.gte_688_48._041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._042_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.gte_688_48._093_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._028_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._036_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._039_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_688_48._027_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48._042_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._043_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_688_48._094_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._029_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._033_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._044_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_688_48._095_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[25] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[24] ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48.B[27] ),
    .D(\efabless_subsystem.compute_controller_i.gte_688_48.B[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._045_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_688_48._096_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[21] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[20] ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48.B[23] ),
    .D(\efabless_subsystem.compute_controller_i.gte_688_48.B[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._046_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_688_48._097_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[17] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[16] ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48.B[19] ),
    .D(\efabless_subsystem.compute_controller_i.gte_688_48.B[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._047_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_688_48._098_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[29] ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48.B[28] ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .D(\efabless_subsystem.compute_controller_i.gte_688_48.B[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._048_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_688_48._099_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48._046_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_688_48._047_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_688_48._048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48._049_ ));
 sky130_fd_sc_hd__a211oi_2 \efabless_subsystem.compute_controller_i.gte_688_48._100_  (.A1(\efabless_subsystem.compute_controller_i.gte_688_48._031_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_688_48._044_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_688_48._045_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_688_48._049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._050_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._000_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._051_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._001_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_700_40._052_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[2] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._000_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._001_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._002_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._053_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._003_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._054_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._004_ ));
 sky130_fd_sc_hd__o211a_2 \efabless_subsystem.compute_controller_i.gte_700_40._055_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[1] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._003_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._004_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40.B[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._005_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_700_40._056_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[2] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._000_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40.B[1] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40._003_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40._005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._006_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._057_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._007_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.gte_700_40._058_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[5] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._008_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._059_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._009_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._060_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._010_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_700_40._061_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._009_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[6] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._010_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._011_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._062_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._012_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_700_40._063_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._012_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._001_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._013_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_700_40._064_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40._008_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40._011_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40._013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._014_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_700_40._065_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._002_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._006_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._015_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_700_40._066_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._010_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[7] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._016_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_700_40._067_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._010_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[7] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._016_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40.B[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._017_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_700_40._068_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._012_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40.B[5] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._018_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_700_40._069_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40._008_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40._011_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40._018_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._019_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._070_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._020_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._071_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._021_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._072_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._022_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_700_40._073_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._023_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._074_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._024_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_700_40._075_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._025_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_700_40._076_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._026_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_700_40._077_  (.A_N(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._027_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.gte_700_40._078_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._024_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._025_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40._026_ ),
    .D1(\efabless_subsystem.compute_controller_i.gte_700_40._027_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._028_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_700_40._079_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._022_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[10] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._023_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40._028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._029_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_700_40._080_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._020_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40._021_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40._029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._030_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.gte_700_40._081_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._015_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._017_ ),
    .A3(\efabless_subsystem.compute_controller_i.gte_700_40._019_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._030_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._031_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_700_40._082_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._020_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40._021_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._032_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.gte_700_40._083_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40.B[9] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._021_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._033_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._084_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._034_ ));
 sky130_fd_sc_hd__or3b_2 \efabless_subsystem.compute_controller_i.gte_700_40._085_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[10] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40._023_ ),
    .C_N(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._035_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_700_40._086_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._034_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[11] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._036_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._087_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._037_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._088_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._038_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_700_40._089_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._037_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[14] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._038_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._039_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_700_40._090_  (.A(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40._040_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_700_40._091_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._024_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40._040_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._041_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_700_40._092_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40._025_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40._026_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40._027_ ),
    .D(\efabless_subsystem.compute_controller_i.gte_700_40._041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._042_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.gte_700_40._093_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._028_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._036_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._039_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_700_40._027_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40._042_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._043_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_700_40._094_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._029_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._033_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._044_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_700_40._095_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[25] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[24] ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40.B[27] ),
    .D(\efabless_subsystem.compute_controller_i.gte_700_40.B[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._045_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_700_40._096_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[21] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[20] ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40.B[23] ),
    .D(\efabless_subsystem.compute_controller_i.gte_700_40.B[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._046_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_700_40._097_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[17] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[16] ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40.B[19] ),
    .D(\efabless_subsystem.compute_controller_i.gte_700_40.B[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._047_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.gte_700_40._098_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[29] ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40.B[28] ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .D(\efabless_subsystem.compute_controller_i.gte_700_40.B[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._048_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.gte_700_40._099_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40._046_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_700_40._047_ ),
    .C(\efabless_subsystem.compute_controller_i.gte_700_40._048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40._049_ ));
 sky130_fd_sc_hd__a211oi_2 \efabless_subsystem.compute_controller_i.gte_700_40._100_  (.A1(\efabless_subsystem.compute_controller_i.gte_700_40._031_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_700_40._044_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_700_40._045_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_700_40._049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.Z ));
 sky130_fd_sc_hd__or3b_2 \efabless_subsystem.compute_controller_i.gte_709_36._1_  (.A(\efabless_subsystem.compute_controller_i.add_163_38.A[0] ),
    .B(\efabless_subsystem.compute_controller_i.add_163_38.A[1] ),
    .C_N(\efabless_subsystem.compute_controller_i._0090_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_709_36._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.gte_709_36._2_  (.A(\efabless_subsystem.compute_controller_i.gte_709_36._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_709_36.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._44_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._00_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._45_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._46_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._02_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_734_31._47_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._48_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._04_ ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.gte_734_31._49_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .B_N(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._05_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.gte_734_31._50_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._04_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._01_ ),
    .B2(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._06_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.gte_734_31._51_  (.A(\efabless_subsystem.compute_controller_i.gte_734_31._04_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .C(\efabless_subsystem.compute_controller_i.gte_734_31._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._07_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_734_31._52_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._00_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._03_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_734_31._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._08_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._53_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._09_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._54_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._55_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._11_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_734_31._56_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._12_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_734_31._57_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._10_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._11_ ),
    .B2(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._13_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_734_31._58_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._14_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._59_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._15_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_734_31._60_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._11_ ),
    .A2(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._15_ ),
    .B2(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._16_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._61_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._17_ ));
 sky130_fd_sc_hd__o2bb2a_2 \efabless_subsystem.compute_controller_i.gte_734_31._62_  (.A1_N(\efabless_subsystem.compute_controller_i.gte_734_31._17_ ),
    .A2_N(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_734_31._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._18_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_734_31._63_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._11_ ),
    .B2(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._19_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_734_31._64_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._12_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._18_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_734_31._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._20_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.gte_734_31._65_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._08_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.gte_734_31._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._21_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._66_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._22_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._67_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._23_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._68_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._24_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._69_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._25_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_734_31._70_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._26_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_734_31._71_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._24_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._25_ ),
    .B2(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._26_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._27_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_734_31._72_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._28_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._73_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._29_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.gte_734_31._74_  (.A(\efabless_subsystem.compute_controller_i.gte_734_31._29_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._30_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._75_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._31_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_734_31._76_  (.A_N(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._32_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_734_31._77_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._31_ ),
    .A2(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._33_ ));
 sky130_fd_sc_hd__o2111a_2 \efabless_subsystem.compute_controller_i.gte_734_31._78_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._28_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._30_ ),
    .D1(\efabless_subsystem.compute_controller_i.gte_734_31._33_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._34_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.compute_controller_i.gte_734_31._79_  (.A(\efabless_subsystem.compute_controller_i.gte_734_31._31_ ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .C(\efabless_subsystem.compute_controller_i.gte_734_31._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._35_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_734_31._80_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._29_ ),
    .B2(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._36_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._81_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._37_ ));
 sky130_fd_sc_hd__a32o_2 \efabless_subsystem.compute_controller_i.gte_734_31._82_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._30_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._33_ ),
    .A3(\efabless_subsystem.compute_controller_i.gte_734_31._36_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._37_ ),
    .B2(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._38_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_734_31._83_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._35_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._38_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._28_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._39_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_734_31._84_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._40_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_734_31._85_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._25_ ),
    .A2(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._40_ ),
    .B2(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._41_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_734_31._86_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_734_31._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31._42_ ));
 sky130_fd_sc_hd__o22ai_2 \efabless_subsystem.compute_controller_i.gte_734_31._87_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._26_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._41_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._42_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_734_31._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_734_31._43_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_734_31._88_  (.A1(\efabless_subsystem.compute_controller_i.gte_734_31._21_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_734_31._34_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_734_31._39_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_734_31._43_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_734_31.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._44_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._00_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._45_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._46_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._02_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_735_31._47_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .B1(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._48_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._04_ ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.gte_735_31._49_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .B_N(\efabless_subsystem.compute_controller_i.gte_286_30.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._05_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.gte_735_31._50_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._04_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._01_ ),
    .B2(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._06_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.gte_735_31._51_  (.A(\efabless_subsystem.compute_controller_i.gte_735_31._04_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .C(\efabless_subsystem.compute_controller_i.gte_735_31._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._07_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_735_31._52_  (.A1(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._00_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._03_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_735_31._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._08_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._53_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._09_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._54_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._55_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._11_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_735_31._56_  (.A_N(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._12_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_735_31._57_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[4] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._10_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._11_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._13_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_735_31._58_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._14_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._59_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._15_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_735_31._60_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._11_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._15_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._16_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._61_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._17_ ));
 sky130_fd_sc_hd__o2bb2a_2 \efabless_subsystem.compute_controller_i.gte_735_31._62_  (.A1_N(\efabless_subsystem.compute_controller_i.gte_735_31._17_ ),
    .A2_N(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_735_31._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._18_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_735_31._63_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._11_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._19_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_735_31._64_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._12_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._18_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_735_31._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._20_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.gte_735_31._65_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._08_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.gte_735_31._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._21_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._66_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._22_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._67_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._23_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._68_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._24_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._69_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._25_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_735_31._70_  (.A_N(\efabless_subsystem.compute_controller_i.acc_cnt_q[15] ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._26_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.gte_735_31._71_  (.A1(\efabless_subsystem.compute_controller_i.gte_286_30.B[13] ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._24_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._25_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[14] ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._26_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._27_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_735_31._72_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._28_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._73_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._29_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.gte_735_31._74_  (.A(\efabless_subsystem.compute_controller_i.gte_735_31._29_ ),
    .B(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._30_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._75_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._31_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.gte_735_31._76_  (.A_N(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._32_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.gte_735_31._77_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._31_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[10] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._33_ ));
 sky130_fd_sc_hd__o2111a_2 \efabless_subsystem.compute_controller_i.gte_735_31._78_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._28_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._30_ ),
    .D1(\efabless_subsystem.compute_controller_i.gte_735_31._33_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._34_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.compute_controller_i.gte_735_31._79_  (.A(\efabless_subsystem.compute_controller_i.gte_735_31._31_ ),
    .B(\efabless_subsystem.compute_controller_i.gte_286_30.B[10] ),
    .C(\efabless_subsystem.compute_controller_i.gte_735_31._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._35_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.gte_735_31._80_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._29_ ),
    .B2(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._36_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._81_  (.A(\efabless_subsystem.compute_controller_i.gte_286_30.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._37_ ));
 sky130_fd_sc_hd__a32o_2 \efabless_subsystem.compute_controller_i.gte_735_31._82_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._30_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._33_ ),
    .A3(\efabless_subsystem.compute_controller_i.gte_735_31._36_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._37_ ),
    .B2(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._38_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.compute_controller_i.gte_735_31._83_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._35_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._38_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._28_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._39_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.gte_735_31._84_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._40_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_735_31._85_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._25_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[14] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._40_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_286_30.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._41_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.gte_735_31._86_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_286_30.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_286_30.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.gte_735_31._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31._42_ ));
 sky130_fd_sc_hd__o22ai_2 \efabless_subsystem.compute_controller_i.gte_735_31._87_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._26_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._41_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._42_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_735_31._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_735_31._43_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.gte_735_31._88_  (.A1(\efabless_subsystem.compute_controller_i.gte_735_31._21_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_735_31._34_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_735_31._39_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_735_31._43_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_735_31.Z ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.lt_156_26._1_  (.A_N(\efabless_subsystem.compute_controller_i.acc_pos_cnt_q ),
    .B(\efabless_subsystem.compute_controller_i._0091_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_156_26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.lt_156_26._2_  (.A(\efabless_subsystem.compute_controller_i.lt_156_26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_156_26.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._48_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._00_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._49_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._01_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.lt_302_35._50_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._00_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._02_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._51_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._52_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._04_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.lt_302_35._53_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._03_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._05_ ));
 sky130_fd_sc_hd__o221a_2 \efabless_subsystem.compute_controller_i.lt_302_35._54_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._00_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._03_ ),
    .B2(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._55_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._07_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.lt_302_35._56_  (.A(\efabless_subsystem.compute_controller_i.lt_302_35._07_ ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._08_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._57_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._09_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._58_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._10_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.lt_302_35._59_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._09_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._11_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._60_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._12_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.lt_302_35._61_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._12_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._13_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.compute_controller_i.lt_302_35._62_  (.A(\efabless_subsystem.compute_controller_i.lt_302_35._08_ ),
    .B(\efabless_subsystem.compute_controller_i.lt_302_35._11_ ),
    .C(\efabless_subsystem.compute_controller_i.lt_302_35._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._14_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.lt_302_35._63_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._02_ ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._06_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._15_ ));
 sky130_fd_sc_hd__o211a_2 \efabless_subsystem.compute_controller_i.lt_302_35._64_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._10_ ),
    .B1(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._16_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.compute_controller_i.lt_302_35._65_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._10_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._17_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.lt_302_35._66_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._12_ ),
    .A2(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._07_ ),
    .B2(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._18_ ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.compute_controller_i.lt_302_35._67_  (.A(\efabless_subsystem.compute_controller_i.lt_302_35._08_ ),
    .B(\efabless_subsystem.compute_controller_i.lt_302_35._11_ ),
    .C(\efabless_subsystem.compute_controller_i.lt_302_35._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._19_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._68_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._20_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._69_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._21_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_controller_i.lt_302_35._70_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[9] ),
    .B(\efabless_subsystem.compute_controller_i.lt_302_35._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._22_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._71_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._23_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._72_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._24_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._73_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._25_ ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.lt_302_35._74_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .B_N(\efabless_subsystem.compute_controller_i.gte_678_56.B[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._26_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.lt_302_35._75_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._25_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._26_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._27_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.lt_302_35._76_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._24_ ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._27_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._28_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._77_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._29_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.lt_302_35._78_  (.A(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.lt_302_35._30_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.lt_302_35._79_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._29_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[10] ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._30_ ),
    .B2(\efabless_subsystem.compute_controller_i.gte_678_56.B[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._31_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.lt_302_35._80_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._20_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._22_ ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._28_ ),
    .D1(\efabless_subsystem.compute_controller_i.lt_302_35._31_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._32_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.lt_302_35._81_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._15_ ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._17_ ),
    .A3(\efabless_subsystem.compute_controller_i.lt_302_35._19_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._32_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._33_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.lt_302_35._82_  (.A_N(\efabless_subsystem.compute_controller_i.gte_678_56.B[15] ),
    .B(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._34_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.lt_302_35._83_  (.A1(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._25_ ),
    .A3(\efabless_subsystem.compute_controller_i.lt_302_35._26_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._34_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._35_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.lt_302_35._84_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._23_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[12] ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[13] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._36_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.lt_302_35._85_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[13] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._24_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._27_ ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._36_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._37_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.lt_302_35._86_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._30_ ),
    .A2(\efabless_subsystem.compute_controller_i.gte_678_56.B[11] ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._29_ ),
    .C1(\efabless_subsystem.compute_controller_i.gte_678_56.B[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._38_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.compute_controller_i.lt_302_35._87_  (.A1(\efabless_subsystem.compute_controller_i.gte_678_56.B[8] ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._20_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[9] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._39_ ));
 sky130_fd_sc_hd__o32a_2 \efabless_subsystem.compute_controller_i.lt_302_35._88_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._22_ ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._31_ ),
    .A3(\efabless_subsystem.compute_controller_i.lt_302_35._39_ ),
    .B1(\efabless_subsystem.compute_controller_i.gte_678_56.B[11] ),
    .B2(\efabless_subsystem.compute_controller_i.lt_302_35._30_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._40_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.lt_302_35._89_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._38_ ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._40_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._28_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._41_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.compute_controller_i.lt_302_35._90_  (.A_N(\efabless_subsystem.compute_controller_i.lt_302_35._35_ ),
    .B(\efabless_subsystem.compute_controller_i.lt_302_35._37_ ),
    .C(\efabless_subsystem.compute_controller_i.lt_302_35._41_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._42_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.lt_302_35._91_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[25] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[24] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[27] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._43_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.lt_302_35._92_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[21] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[20] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[23] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._44_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.lt_302_35._93_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[17] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[16] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[19] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._45_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.lt_302_35._94_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[29] ),
    .B(\efabless_subsystem.compute_controller_i.gte_678_56.B[28] ),
    .C(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .D(\efabless_subsystem.compute_controller_i.gte_678_56.B[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._46_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.lt_302_35._95_  (.A(\efabless_subsystem.compute_controller_i.lt_302_35._44_ ),
    .B(\efabless_subsystem.compute_controller_i.lt_302_35._45_ ),
    .C(\efabless_subsystem.compute_controller_i.lt_302_35._46_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35._47_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.lt_302_35._96_  (.A1(\efabless_subsystem.compute_controller_i.lt_302_35._33_ ),
    .A2(\efabless_subsystem.compute_controller_i.lt_302_35._42_ ),
    .B1(\efabless_subsystem.compute_controller_i.lt_302_35._43_ ),
    .C1(\efabless_subsystem.compute_controller_i.lt_302_35._47_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.lt_302_35.Z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[15] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[15] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[6] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[6] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[5] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[5] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[4] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[3] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[2] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[1] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[0] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[14] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[14] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[13] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[13] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[12] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[12] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[11] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[11] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[10] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[10] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[9] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[9] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[8] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[8] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_185_30.Z[7] ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_cnt_d[7] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[15] ),
    .A1(\efabless_subsystem.compute_controller_i._0364_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g10._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[6] ),
    .A1(\efabless_subsystem.compute_controller_i._0355_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g10._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g10.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g11._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[5] ),
    .A1(\efabless_subsystem.compute_controller_i._0354_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g11._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g11.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g12._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[4] ),
    .A1(\efabless_subsystem.compute_controller_i._0353_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g12._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g12.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g13._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0352_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g13._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g13.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g14._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0351_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g14._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g14.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g15._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0350_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g15._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g15.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g16._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0349_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g16._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g16.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[14] ),
    .A1(\efabless_subsystem.compute_controller_i._0363_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[13] ),
    .A1(\efabless_subsystem.compute_controller_i._0362_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[12] ),
    .A1(\efabless_subsystem.compute_controller_i._0361_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g5._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[11] ),
    .A1(\efabless_subsystem.compute_controller_i._0360_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g5._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g5.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g6._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[10] ),
    .A1(\efabless_subsystem.compute_controller_i._0359_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g6._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g6.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g7._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[9] ),
    .A1(\efabless_subsystem.compute_controller_i._0358_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g7._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g7.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g8._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[8] ),
    .A1(\efabless_subsystem.compute_controller_i._0357_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g8._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g8.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g9._1_  (.A0(\efabless_subsystem.compute_controller_i.acc_cnt_q[7] ),
    .A1(\efabless_subsystem.compute_controller_i._0356_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g9._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_190_15.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_cnt_d_184_9.g9.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0365_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_pos_cnt_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_156_26.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0366_ ),
    .A1(\efabless_subsystem.compute_controller_i.add_157_42.Z ),
    .S(\efabless_subsystem.compute_controller_i.lt_156_26.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_156_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_156_26.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_156_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._3_  (.A1(\efabless_subsystem.compute_controller_i._0367_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[3] ),
    .B1(\efabless_subsystem.compute_controller_i._0092_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._0_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._4_  (.A1(\efabless_subsystem.compute_controller_i._0368_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[1] ),
    .B1(\efabless_subsystem.compute_controller_i._0369_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._1_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._5_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._0_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._6_  (.A(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2].d ),
    .A1(\efabless_subsystem.compute_controller_i._0372_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_d[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1].d ),
    .A1(\efabless_subsystem.compute_controller_i._0371_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_654_22.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_d[1] ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._3_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data1 ),
    .A2(\efabless_subsystem.compute_controller_i._0374_ ),
    .A3(\efabless_subsystem.compute_controller_i._0376_ ),
    .S0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._0_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._4_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data2 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data3 ),
    .A2(\efabless_subsystem.compute_controller_i._0379_ ),
    .A3(\efabless_subsystem.compute_controller_i._0382_ ),
    .S0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._1_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._5_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._0_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._1_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._6_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[2].d ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._3_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data1 ),
    .A2(\efabless_subsystem.compute_controller_i._0373_ ),
    .A3(\efabless_subsystem.compute_controller_i._0375_ ),
    .S0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._0_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._4_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data2 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data3 ),
    .A2(\efabless_subsystem.compute_controller_i._0378_ ),
    .A3(\efabless_subsystem.compute_controller_i._0381_ ),
    .S0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._1_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._5_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._0_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._1_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._6_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[1].d ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._3_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data1 ),
    .A2(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data4 ),
    .A3(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data5 ),
    .S0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._0_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._4_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data2 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data3 ),
    .A2(\efabless_subsystem.compute_controller_i._0377_ ),
    .A3(\efabless_subsystem.compute_controller_i._0380_ ),
    .S0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._1_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._5_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._0_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._1_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._6_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0384_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0383_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0093_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0095_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0385_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0094_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0096_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_688_48.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0387_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_688_48.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0386_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_688_48.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_688_48.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_683_39.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0389_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0097_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0388_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_694_44.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_678_21.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0390_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0099_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0098_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_700_40.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_700_40.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_672_66.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0101_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0391_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0100_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_710_18.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0103_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g1.data3 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0392_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g2.data3 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.arr_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0102_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_720_66.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data3 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0104_ ),
    .A1(\efabless_subsystem.compute_controller_i._0393_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data4 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_749_18.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0105_ ),
    .A1(\efabless_subsystem.compute_controller_i._0394_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_735_18.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_749_18.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_749_18.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_749_18.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_659_15.g3.data5 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0396_ ),
    .A1(\efabless_subsystem.compute_controller_i.add_163_38.Z[1] ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_d[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g2._1_  (.A0(\efabless_subsystem.compute_controller_i._0395_ ),
    .A1(\efabless_subsystem.compute_controller_i.add_163_38.Z[0] ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_pos_cnt_d_153_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_aux_pos_cnt_d_153_6.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.aux_pos_cnt_d[0] ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._08_  (.A1(\efabless_subsystem.compute_controller_i._0423_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[9] ),
    .B1(\efabless_subsystem.compute_controller_i._0419_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._00_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._09_  (.A1(\efabless_subsystem.compute_controller_i._0408_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[10] ),
    .B1(\efabless_subsystem.compute_controller_i._0430_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._01_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._10_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._00_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._02_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._11_  (.A1(\efabless_subsystem.compute_controller_i._0443_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[4] ),
    .B1(\efabless_subsystem.compute_controller_i._0413_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._03_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._12_  (.A1(\efabless_subsystem.compute_controller_i._0402_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[11] ),
    .B1(\efabless_subsystem.compute_controller_i._0450_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[2] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._04_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._13_  (.A1(\efabless_subsystem.compute_controller_i._0111_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[8] ),
    .B1(\efabless_subsystem.compute_controller_i._0435_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._05_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._14_  (.A1(\efabless_subsystem.compute_controller_i._0439_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[5] ),
    .B1(\efabless_subsystem.compute_controller_i._0447_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[3] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._06_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._15_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._02_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._04_ ),
    .C(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._16_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g1._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_arr_fsm_state_d_663_21.ctl ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._08_  (.A1(\efabless_subsystem.compute_controller_i._0108_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[9] ),
    .B1(\efabless_subsystem.compute_controller_i._0418_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._00_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._09_  (.A1(\efabless_subsystem.compute_controller_i._0407_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[10] ),
    .B1(\efabless_subsystem.compute_controller_i._0113_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._01_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._10_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._00_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._02_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._11_  (.A1(\efabless_subsystem.compute_controller_i._0118_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[4] ),
    .B1(\efabless_subsystem.compute_controller_i._0412_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._03_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._12_  (.A1(\efabless_subsystem.compute_controller_i._0401_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[11] ),
    .B1(\efabless_subsystem.compute_controller_i._0123_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[2] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._04_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._13_  (.A1(\efabless_subsystem.compute_controller_i._0110_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[8] ),
    .B1(\efabless_subsystem.compute_controller_i._0114_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._05_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._14_  (.A1(\efabless_subsystem.compute_controller_i._0116_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[5] ),
    .B1(\efabless_subsystem.compute_controller_i._0120_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[3] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._06_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._15_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._02_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._04_ ),
    .C(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._16_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g2.z ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._08_  (.A1(\efabless_subsystem.compute_controller_i._0420_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[9] ),
    .B1(\efabless_subsystem.compute_controller_i._0414_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._00_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._09_  (.A1(\efabless_subsystem.compute_controller_i._0403_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[10] ),
    .B1(\efabless_subsystem.compute_controller_i._0427_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._01_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._10_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._00_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._02_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._11_  (.A1(\efabless_subsystem.compute_controller_i._0440_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[4] ),
    .B1(\efabless_subsystem.compute_controller_i._0106_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._03_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._12_  (.A1(\efabless_subsystem.compute_controller_i._0397_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[11] ),
    .B1(\efabless_subsystem.compute_controller_i._0448_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[2] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._04_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._13_  (.A1(\efabless_subsystem.compute_controller_i._0424_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[8] ),
    .B1(\efabless_subsystem.compute_controller_i._0431_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._05_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._14_  (.A1(\efabless_subsystem.compute_controller_i._0436_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[5] ),
    .B1(\efabless_subsystem.compute_controller_i._0444_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_375_11.out_0[3] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._06_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._15_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._02_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._04_ ),
    .C(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._16_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_array_start_375_11.g6._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_done ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._3_  (.A1(\efabless_subsystem.compute_controller_i._0124_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[5] ),
    .B1(\efabless_subsystem.compute_controller_i._0455_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._0_ ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._4_  (.A1(\efabless_subsystem.compute_controller_i._0452_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[6] ),
    .B1(\efabless_subsystem.compute_controller_i._0457_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._1_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._5_  (.A1(\efabless_subsystem.compute_controller_i._0126_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[2] ),
    .B1(\efabless_subsystem.compute_controller_i._0458_ ),
    .B2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[1] ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._2_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._6_  (.A1(\efabless_subsystem.compute_controller_i._0460_ ),
    .A2(\efabless_subsystem.compute_controller_i.ctl_775_11.out_0[0] ),
    .B1(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._0_ ),
    .C1(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1.z ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._15_  (.A0(\efabless_subsystem.compute_controller_i._0464_ ),
    .A1(\efabless_subsystem.compute_controller_i._0468_ ),
    .A2(\efabless_subsystem.compute_controller_i._0480_ ),
    .A3(\efabless_subsystem.compute_controller_i._0484_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._16_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._17_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data7 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._02_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._18_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i._0487_ ),
    .B1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._03_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._19_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._03_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._20_  (.A(\efabless_subsystem.compute_controller_i._0486_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._21_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._06_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._22_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._05_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._07_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._23_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._08_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._24_  (.A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._04_ ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._07_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._09_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._25_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data8 ),
    .A1(\efabless_subsystem.compute_controller_i._0488_ ),
    .A2(\efabless_subsystem.compute_controller_i._0472_ ),
    .A3(\efabless_subsystem.compute_controller_i._0476_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._26_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._11_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._27_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data1 ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data4 ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data5 ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._12_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._28_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._13_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._29_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._13_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._14_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._30_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._09_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[3].d ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._15_  (.A0(\efabless_subsystem.compute_controller_i._0463_ ),
    .A1(\efabless_subsystem.compute_controller_i._0467_ ),
    .A2(\efabless_subsystem.compute_controller_i._0479_ ),
    .A3(\efabless_subsystem.compute_controller_i._0483_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._16_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._17_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data7 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._02_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._18_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i._0131_ ),
    .B1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._03_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._19_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._03_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._20_  (.A(\efabless_subsystem.compute_controller_i._0128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._21_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._06_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._22_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._05_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._07_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._23_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._08_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._24_  (.A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._04_ ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._07_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._09_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._25_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data8 ),
    .A1(\efabless_subsystem.compute_controller_i._0134_ ),
    .A2(\efabless_subsystem.compute_controller_i._0471_ ),
    .A3(\efabless_subsystem.compute_controller_i._0475_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._26_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._11_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._27_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data1 ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data4 ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data5 ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._12_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._28_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._13_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._29_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._13_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._14_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._30_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._09_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[2].d ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._15_  (.A0(\efabless_subsystem.compute_controller_i._0462_ ),
    .A1(\efabless_subsystem.compute_controller_i._0466_ ),
    .A2(\efabless_subsystem.compute_controller_i._0478_ ),
    .A3(\efabless_subsystem.compute_controller_i._0482_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._16_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._17_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data7 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._02_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._18_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i._0130_ ),
    .B1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._03_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._19_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._03_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._20_  (.A(\efabless_subsystem.compute_controller_i._0485_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._21_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._06_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._22_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._05_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._07_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._23_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._08_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._24_  (.A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._04_ ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._07_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._09_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._25_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data8 ),
    .A1(\efabless_subsystem.compute_controller_i._0133_ ),
    .A2(\efabless_subsystem.compute_controller_i._0470_ ),
    .A3(\efabless_subsystem.compute_controller_i._0474_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._26_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._11_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._27_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data1 ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data4 ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data5 ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._12_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._28_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._13_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._29_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._13_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._14_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._30_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._09_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[1].d ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._15_  (.A0(\efabless_subsystem.compute_controller_i._0461_ ),
    .A1(\efabless_subsystem.compute_controller_i._0465_ ),
    .A2(\efabless_subsystem.compute_controller_i._0477_ ),
    .A3(\efabless_subsystem.compute_controller_i._0481_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._16_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._17_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data7 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._02_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._18_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i._0129_ ),
    .B1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._03_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._19_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._03_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._20_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data3 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._21_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._06_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._22_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._05_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._06_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .D1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._07_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._23_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._08_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._24_  (.A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._01_ ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._04_ ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._07_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._09_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._25_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data8 ),
    .A1(\efabless_subsystem.compute_controller_i._0132_ ),
    .A2(\efabless_subsystem.compute_controller_i._0469_ ),
    .A3(\efabless_subsystem.compute_controller_i._0473_ ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._10_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._26_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._11_ ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._27_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data1 ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data4 ),
    .A3(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data5 ),
    .S0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .S1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._12_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._28_  (.A(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._13_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._29_  (.A1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A2(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._13_ ),
    .C1(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._14_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._30_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._09_ ),
    .B(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0491_ ),
    .S(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0490_ ),
    .S(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0489_ ),
    .S(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0135_ ),
    .S(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_248_21.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0494_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_255_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0493_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_255_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0136_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_255_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0492_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_255_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_255_34.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0496_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0495_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0138_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0137_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_262_34.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_269_32.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0139_ ),
    .A1(\efabless_subsystem.compute_controller_i._0497_ ),
    .S(\efabless_subsystem.compute_controller_i.gt_269_32.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_269_32.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_269_32.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_269_32.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data3 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0499_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data4 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0141_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data4 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0498_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data4 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0140_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_278_34.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data4 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0501_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data5 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0143_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data5 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0142_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data5 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0500_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data5 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1.data1 ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data7 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2.data1 ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data7 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3.data1 ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data7 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4.data1 ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data7 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0144_ ),
    .S(\efabless_subsystem.compute_controller_i.lt_302_35.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0504_ ),
    .S(\efabless_subsystem.compute_controller_i.lt_302_35.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0503_ ),
    .S(\efabless_subsystem.compute_controller_i.lt_302_35.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0502_ ),
    .S(\efabless_subsystem.compute_controller_i.lt_302_35.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_299_34.g4.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0506_ ),
    .A1(\efabless_subsystem.compute_controller_i._0148_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_734_31.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g2._1_  (.A0(\efabless_subsystem.compute_controller_i._0146_ ),
    .A1(\efabless_subsystem.compute_controller_i._0508_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_734_31.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g3._1_  (.A0(\efabless_subsystem.compute_controller_i._0505_ ),
    .A1(\efabless_subsystem.compute_controller_i._0147_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_734_31.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g4._1_  (.A0(\efabless_subsystem.compute_controller_i._0145_ ),
    .A1(\efabless_subsystem.compute_controller_i._0507_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_734_31.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_308_39.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_302_35.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0150_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g1.data8 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0510_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g2.data8 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0509_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g3.data8 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0149_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_244_15.g4.data8 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0511_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0151_ ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[1] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3.data1 ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.context_fsm_state_q[0] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4.data1 ),
    .S(\efabless_subsystem.compute_controller_i.gte_262_34.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_324_17.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0512_ ),
    .A1(\efabless_subsystem.compute_controller_i._0153_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g2._1_  (.A0(\efabless_subsystem.compute_controller_i._0152_ ),
    .A1(\efabless_subsystem.compute_controller_i._0513_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_286_17.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_333_21.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_context_fsm_state_d_329_43.g4.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[15] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[15] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[6] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[6] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[5] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[5] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[4] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[3] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[2] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[1] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[0] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[14] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[14] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[13] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[13] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[12] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[12] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[11] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[11] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[10] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[10] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[9] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[9] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[8] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[8] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9.data0 ),
    .A1(\efabless_subsystem.compute_controller_i.add_200_30.Z[7] ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.ctx_cnt_d[7] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[15] ),
    .A1(\efabless_subsystem.compute_controller_i._0529_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g10._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[6] ),
    .A1(\efabless_subsystem.compute_controller_i._0520_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g10._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g10.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g11._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[5] ),
    .A1(\efabless_subsystem.compute_controller_i._0519_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g11._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g11.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g12._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[4] ),
    .A1(\efabless_subsystem.compute_controller_i._0518_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g12._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g12.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g13._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[3] ),
    .A1(\efabless_subsystem.compute_controller_i._0517_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g13._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g13.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g14._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[2] ),
    .A1(\efabless_subsystem.compute_controller_i._0516_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g14._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g14.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g15._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0515_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g15._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g15.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g16._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0514_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g16._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g16.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[14] ),
    .A1(\efabless_subsystem.compute_controller_i._0528_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[13] ),
    .A1(\efabless_subsystem.compute_controller_i._0527_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[12] ),
    .A1(\efabless_subsystem.compute_controller_i._0526_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g5._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[11] ),
    .A1(\efabless_subsystem.compute_controller_i._0525_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g5._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g5.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g6._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[10] ),
    .A1(\efabless_subsystem.compute_controller_i._0524_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g6._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g6.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g7._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[9] ),
    .A1(\efabless_subsystem.compute_controller_i._0523_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g7._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g7.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g8._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[8] ),
    .A1(\efabless_subsystem.compute_controller_i._0522_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g8._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g8.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g9._1_  (.A0(\efabless_subsystem.compute_controller_i.add_200_30.A[7] ),
    .A1(\efabless_subsystem.compute_controller_i._0521_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g9._2_  (.A(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_203_38.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_ctx_cnt_d_198_6.g9.data0 ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0154_ ),
    .A2(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.data2 ),
    .A3(\efabless_subsystem.compute_controller_i._0532_ ),
    .S0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .S1(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.z ));
 sky130_fd_sc_hd__mux4_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.data0 ),
    .A1(\efabless_subsystem.compute_controller_i._0530_ ),
    .A2(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.data2 ),
    .A3(\efabless_subsystem.compute_controller_i._0531_ ),
    .S0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .S1(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0533_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .A1(\efabless_subsystem.compute_controller_i._0155_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_557_53.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .A1(\efabless_subsystem.compute_controller_i._0534_ ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2.data1 ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_edge ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.data2 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0535_ ),
    .A1(\efabless_subsystem.compute_controller_i._0156_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_575_57.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_571_21.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0551_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10._1_  (.A0(\efabless_subsystem.compute_controller_i._0542_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11._1_  (.A0(\efabless_subsystem.compute_controller_i._0541_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12._1_  (.A0(\efabless_subsystem.compute_controller_i._0540_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13._1_  (.A0(\efabless_subsystem.compute_controller_i._0539_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14._1_  (.A0(\efabless_subsystem.compute_controller_i._0538_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15._1_  (.A0(\efabless_subsystem.compute_controller_i._0537_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16._1_  (.A0(\efabless_subsystem.compute_controller_i._0536_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2._1_  (.A0(\efabless_subsystem.compute_controller_i._0550_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3._1_  (.A0(\efabless_subsystem.compute_controller_i._0549_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4._1_  (.A0(\efabless_subsystem.compute_controller_i._0548_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5._1_  (.A0(\efabless_subsystem.compute_controller_i._0547_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6._1_  (.A0(\efabless_subsystem.compute_controller_i._0546_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7._1_  (.A0(\efabless_subsystem.compute_controller_i._0545_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8._1_  (.A0(\efabless_subsystem.compute_controller_i._0544_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9._1_  (.A0(\efabless_subsystem.compute_controller_i._0543_ ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9.data1 ),
    .S(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g1._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[15] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g10._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[6] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g10._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g11._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[5] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g11._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g12._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[4] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g12._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g13._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[3] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g13._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g14._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[2] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g14._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g15._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[1] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g15._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g16._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[0] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g16._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g2._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[14] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g2._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g3._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[13] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g3._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g4._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[12] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g4._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g5._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[11] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g5._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g6._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[10] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g6._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g7._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[9] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g7._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g8._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[8] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g8._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g9._1_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .A1(\efabless_subsystem.compute_controller_i.add_175_34.Z[7] ),
    .S(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g9._2_  (.A(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_174_13.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1._1_  (.A0(\efabless_subsystem.compute_controller_i._0552_ ),
    .A1(\efabless_subsystem.compute_controller_i.add_143_38.Z ),
    .S(\efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1._2_  (.A(\efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1.z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g2.z ),
    .S(\efabless_subsystem.compute_controller_i._0157_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0554_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0555_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_psm_fsm_state_d_553_15.g1.z ),
    .S(\efabless_subsystem.compute_controller_i._0158_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0556_ ),
    .S(\efabless_subsystem.compute_controller_i.arr_fsm_state_q_reg[0].srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.ctl_psm_fsm_state_q_603_11.in_0[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.psm_fsm_state_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0557_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g16.z ),
    .S(\efabless_subsystem.compute_controller_i._0159_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0558_ ),
    .S(\efabless_subsystem.compute_controller_i._0559_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[0] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0560_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g6.z ),
    .S(\efabless_subsystem.compute_controller_i._0160_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0561_ ),
    .S(\efabless_subsystem.compute_controller_i._0562_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[10] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g5.z ),
    .S(\efabless_subsystem.compute_controller_i._0161_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0564_ ),
    .S(\efabless_subsystem.compute_controller_i._0565_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[11] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0566_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g4.z ),
    .S(\efabless_subsystem.compute_controller_i._0162_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0567_ ),
    .S(\efabless_subsystem.compute_controller_i._0568_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[12] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0569_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g3.z ),
    .S(\efabless_subsystem.compute_controller_i._0163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0570_ ),
    .S(\efabless_subsystem.compute_controller_i._0571_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[13] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[13]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0572_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g2.z ),
    .S(\efabless_subsystem.compute_controller_i._0164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0573_ ),
    .S(\efabless_subsystem.compute_controller_i._0574_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[14] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[14]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0575_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g1.z ),
    .S(\efabless_subsystem.compute_controller_i._0165_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0576_ ),
    .S(\efabless_subsystem.compute_controller_i._0577_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[15] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[15]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0578_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g15.z ),
    .S(\efabless_subsystem.compute_controller_i._0166_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0579_ ),
    .S(\efabless_subsystem.compute_controller_i._0580_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[1] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0581_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g14.z ),
    .S(\efabless_subsystem.compute_controller_i._0167_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0582_ ),
    .S(\efabless_subsystem.compute_controller_i._0583_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[2] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0584_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g13.z ),
    .S(\efabless_subsystem.compute_controller_i._0168_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0585_ ),
    .S(\efabless_subsystem.compute_controller_i._0586_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[3] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0587_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g12.z ),
    .S(\efabless_subsystem.compute_controller_i._0169_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0588_ ),
    .S(\efabless_subsystem.compute_controller_i._0589_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[4] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0590_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g11.z ),
    .S(\efabless_subsystem.compute_controller_i._0170_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0591_ ),
    .S(\efabless_subsystem.compute_controller_i._0592_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[5] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0593_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g10.z ),
    .S(\efabless_subsystem.compute_controller_i._0171_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0594_ ),
    .S(\efabless_subsystem.compute_controller_i._0595_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[6] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0596_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g9.z ),
    .S(\efabless_subsystem.compute_controller_i._0172_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0597_ ),
    .S(\efabless_subsystem.compute_controller_i._0598_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[7] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0599_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g8.z ),
    .S(\efabless_subsystem.compute_controller_i._0173_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0600_ ),
    .S(\efabless_subsystem.compute_controller_i._0601_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[8] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._08_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0602_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .A1(\efabless_subsystem.compute_controller_i.mux_red_cnt_d_173_26.g7.z ),
    .S(\efabless_subsystem.compute_controller_i._0174_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._10_  (.A0(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0603_ ),
    .S(\efabless_subsystem.compute_controller_i._0604_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._11_  (.A(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_175_34.A[9] ),
    .Q_N(\efabless_subsystem.compute_controller_i.red_cnt_q_reg[9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_controller_i.acc_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_controller_i._0605_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_controller_i.add_143_38.A ),
    .A1(\efabless_subsystem.compute_controller_i.mux_startup_cnt_d_142_29.g1.z ),
    .S(\efabless_subsystem.compute_controller_i._0175_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_controller_i._0606_ ),
    .S(\efabless_subsystem.compute_controller_i._0607_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.add_143_38.A ),
    .Q_N(\efabless_subsystem.compute_controller_i.startup_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__or3b_2 \efabless_subsystem.compute_controller_i.sub_302_49._22_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[1] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .C_N(\efabless_subsystem.compute_controller_i._0176_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.sub_302_49._23_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.sub_302_49._24_  (.A(\efabless_subsystem.compute_controller_i._0176_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_302_49._02_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_302_49._25_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_302_49._03_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_302_49._26_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._01_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[1] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._27_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[2] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._28_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._04_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_302_49._29_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._01_ ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_302_49._05_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_302_49._30_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._04_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._31_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[4] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._32_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._06_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_302_49._33_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._04_ ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_302_49._07_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_302_49._34_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._06_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[5] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._35_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[6] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_302_49._36_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .D(\efabless_subsystem.compute_controller_i.sub_302_49._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._08_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_302_49._37_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .D(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._09_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_302_49._38_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._01_ ),
    .D(\efabless_subsystem.compute_controller_i.sub_302_49._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.sub_302_49._39_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_302_49._40_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._08_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[7] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._41_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[8] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._42_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._12_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_302_49._43_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_302_49._13_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_302_49._44_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._12_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[9] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._45_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._14_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.sub_302_49._46_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._15_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_302_49._47_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._12_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_302_49._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[10] ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.sub_302_49._48_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._16_ ));
 sky130_fd_sc_hd__a2bb2o_2 \efabless_subsystem.compute_controller_i.sub_302_49._49_  (.A1_N(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .A2_N(\efabless_subsystem.compute_controller_i.sub_302_49._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_302_49._15_ ),
    .B2(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[11] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._50_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._17_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_302_49._51_  (.A1(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_302_49._18_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_302_49._52_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._17_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[12] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_302_49._53_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .D(\efabless_subsystem.compute_controller_i.sub_302_49._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._19_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_302_49._54_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._17_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_302_49._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[13] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._55_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .B(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .C(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._20_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_302_49._56_  (.A(\efabless_subsystem.compute_controller_i.sub_302_49._11_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._16_ ),
    .C(\efabless_subsystem.compute_controller_i.sub_302_49._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_302_49._21_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_302_49._57_  (.A1(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_302_49._19_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_302_49._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[14] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._58_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[15] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._59_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .B(\efabless_subsystem.compute_controller_i._0176_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[0] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.sub_302_49._60_  (.A(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .B(\efabless_subsystem.compute_controller_i.sub_302_49._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._61_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._62_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._63_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._64_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._65_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._66_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._67_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._68_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._69_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._70_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._71_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._72_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._73_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._74_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_302_49._75_  (.A(\efabless_subsystem.compute_controller_i.gte_678_56.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_678_56.B[30] ));
 sky130_fd_sc_hd__nand2b_2 \efabless_subsystem.compute_controller_i.sub_688_68._25_  (.A_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .B(\efabless_subsystem.compute_controller_i._0608_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._00_ ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.sub_688_68._26_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ),
    .B_N(\efabless_subsystem.compute_controller_i._0177_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.sub_688_68._27_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._02_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.sub_688_68._28_  (.A_N(\efabless_subsystem.compute_controller_i._0177_ ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._29_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._02_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._04_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._30_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._00_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[1] ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.sub_688_68._31_  (.A1(\efabless_subsystem.compute_controller_i.sub_688_68._00_ ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._01_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_688_68._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._05_ ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._32_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[2] ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.sub_688_68._33_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._06_ ));
 sky130_fd_sc_hd__a211o_2 \efabless_subsystem.compute_controller_i.sub_688_68._34_  (.A1(\efabless_subsystem.compute_controller_i.sub_688_68._00_ ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._01_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_688_68._03_ ),
    .C1(\efabless_subsystem.compute_controller_i.sub_688_68._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._07_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_688_68._35_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._05_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._08_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_688_68._36_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._07_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._37_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[4] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_688_68._38_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.sub_688_68._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._09_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_688_68._39_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._07_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._10_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_688_68._40_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._09_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[5] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._41_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[6] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_688_68._42_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .D(\efabless_subsystem.compute_controller_i.sub_688_68._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._11_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_688_68._43_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._12_ ));
 sky130_fd_sc_hd__a2111o_2 \efabless_subsystem.compute_controller_i.sub_688_68._44_  (.A1(\efabless_subsystem.compute_controller_i.sub_688_68._00_ ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._01_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_688_68._03_ ),
    .C1(\efabless_subsystem.compute_controller_i.sub_688_68._06_ ),
    .D1(\efabless_subsystem.compute_controller_i.sub_688_68._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_688_68._45_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._11_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[7] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._46_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[8] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_688_68._47_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._14_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_688_68._48_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._15_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_688_68._49_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._14_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[9] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_688_68._50_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .D(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._16_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_688_68._51_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._14_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_688_68._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[10] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_688_68._52_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._17_ ));
 sky130_fd_sc_hd__a2bb2o_2 \efabless_subsystem.compute_controller_i.sub_688_68._53_  (.A1_N(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .A2_N(\efabless_subsystem.compute_controller_i.sub_688_68._17_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_688_68._16_ ),
    .B2(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[11] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_688_68._54_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .C(\efabless_subsystem.compute_controller_i.sub_688_68._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._18_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_688_68._55_  (.A1(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._17_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._19_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_688_68._56_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._18_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[12] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_688_68._57_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .C(\efabless_subsystem.compute_controller_i.sub_688_68._17_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._20_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.sub_688_68._58_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._21_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_688_68._59_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._18_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_688_68._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[13] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.compute_controller_i.sub_688_68._60_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._13_ ),
    .C(\efabless_subsystem.compute_controller_i.sub_688_68._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_688_68._22_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_controller_i.sub_688_68._61_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_688_68._21_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_688_68._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[14] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.sub_688_68._62_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[15] ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_controller_i.sub_688_68._63_  (.A(\efabless_subsystem.compute_controller_i._0608_ ),
    .B_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._23_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_688_68._64_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._00_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._23_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_688_48.B[0] ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_controller_i.sub_688_68._65_  (.A_N(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ),
    .B(\efabless_subsystem.compute_controller_i.sub_688_68._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_688_68._24_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.sub_688_68._66_  (.A(\efabless_subsystem.compute_controller_i.sub_688_68._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._67_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._68_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._69_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._70_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._71_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._72_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._73_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._74_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._75_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._76_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._77_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._78_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._79_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._80_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_688_68._81_  (.A(\efabless_subsystem.compute_controller_i.gte_688_48.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_688_48.B[30] ));
 sky130_fd_sc_hd__or3b_2 \efabless_subsystem.compute_controller_i.sub_700_60._22_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .C_N(\efabless_subsystem.compute_controller_i._0178_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.sub_700_60._23_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_controller_i.sub_700_60._24_  (.A(\efabless_subsystem.compute_controller_i._0178_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_700_60._02_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_700_60._25_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._02_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_700_60._03_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_700_60._26_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._01_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[1] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._27_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[2] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._28_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._04_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_700_60._29_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._01_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_700_60._05_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_700_60._30_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._04_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._31_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[4] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._32_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._06_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_700_60._33_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._04_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_700_60._07_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_700_60._34_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._06_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[5] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._35_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[6] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_700_60._36_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .D(\efabless_subsystem.compute_controller_i.sub_700_60._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._08_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_700_60._37_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[4] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[5] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[6] ),
    .D(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._09_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_700_60._38_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[2] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[3] ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._01_ ),
    .D(\efabless_subsystem.compute_controller_i.sub_700_60._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_controller_i.sub_700_60._39_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_700_60._40_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[7] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._08_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[7] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._41_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[8] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._42_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._12_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_700_60._43_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_700_60._13_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_700_60._44_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._12_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[9] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._45_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[8] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[9] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._14_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.sub_700_60._46_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._15_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_700_60._47_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[10] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._12_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_700_60._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[10] ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_controller_i.sub_700_60._48_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._16_ ));
 sky130_fd_sc_hd__a2bb2o_2 \efabless_subsystem.compute_controller_i.sub_700_60._49_  (.A1_N(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .A2_N(\efabless_subsystem.compute_controller_i.sub_700_60._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.sub_700_60._15_ ),
    .B2(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[11] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._50_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._17_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.compute_controller_i.sub_700_60._51_  (.A1(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._16_ ),
    .B1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.sub_700_60._18_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_controller_i.sub_700_60._52_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._17_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[12] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.compute_controller_i.sub_700_60._53_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .D(\efabless_subsystem.compute_controller_i.sub_700_60._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._19_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_700_60._54_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._17_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_700_60._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[13] ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._55_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[12] ),
    .B(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[13] ),
    .C(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._20_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.compute_controller_i.sub_700_60._56_  (.A(\efabless_subsystem.compute_controller_i.sub_700_60._11_ ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._16_ ),
    .C(\efabless_subsystem.compute_controller_i.sub_700_60._20_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.sub_700_60._21_ ));
 sky130_fd_sc_hd__a21bo_2 \efabless_subsystem.compute_controller_i.sub_700_60._57_  (.A1(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[14] ),
    .A2(\efabless_subsystem.compute_controller_i.sub_700_60._19_ ),
    .B1_N(\efabless_subsystem.compute_controller_i.sub_700_60._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[14] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._58_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[15] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._59_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[0] ),
    .B(\efabless_subsystem.compute_controller_i._0178_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[0] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.compute_controller_i.sub_700_60._60_  (.A(\efabless_subsystem.compute_controller_i.arr_red_cycles_q[15] ),
    .B(\efabless_subsystem.compute_controller_i.sub_700_60._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._61_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._62_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._63_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._64_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._65_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._66_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._67_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._68_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._69_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._70_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._71_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._72_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._73_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._74_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_controller_i.sub_700_60._75_  (.A(\efabless_subsystem.compute_controller_i.gte_700_40.B[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.gte_700_40.B[30] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_core_i._2_  (.A(\efabless_subsystem.compute_core_i.shftsgn_reg_valid ),
    .B(\efabless_subsystem.compute_core_i.weight_reg_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i._3_  (.A(\efabless_subsystem.compute_core_i._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.mux_152_27.g1.data1 ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_core_i._4_  (.A(\efabless_subsystem.compute_core_i.shftsgn_reg_valid ),
    .B(\efabless_subsystem.compute_core_i.fmap_reg_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i._1_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i._5_  (.A(\efabless_subsystem.compute_core_i._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.mux_152_27.g1.data0 ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.compute_core_i.array_accumulator_i._653_  (.A(\efabless_subsystem.compute_controller_i.mux_cmbsop_o_pipeline_ready_775_11.g1.z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.array_acc_ready ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._143_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_reg_q_reg[0][0].aclr ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._144_  (.A(\efabless_subsystem.compute_core_i.array_acc_ready ),
    .B_N(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._000_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._145_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._000_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_ready_i ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._148_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._002_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._149_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._002_ ),
    .B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_ready_i ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._003_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._150_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._285_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._137_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._286_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._138_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._287_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._139_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._288_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._140_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._289_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._141_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._290_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._142_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._07_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_reg_q_reg[0][0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._08_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._137_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._09_  (.A0(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid ),
    .A1(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0].d ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_ready_i ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._10_  (.A0(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._138_ ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._11_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid ),
    .Q_N(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._07_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_reg_q_reg[0][0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._08_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._140_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._09_  (.A0(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .A1(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_ready_i ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._10_  (.A0(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._141_ ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i._142_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._11_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.i_arr_data_valid ),
    .Q_N(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.ifmap_regs_i._07_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0].aclr ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.ifmap_regs_i._08_  (.A0(\efabless_subsystem.compute_core_i.fmap_reg_valid ),
    .A1(\efabless_subsystem.compute_core_i.i_fmap_valid ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.ifmap_regs_i._09_  (.A(\efabless_subsystem.compute_core_i.ifmap_regs_i._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_d ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_core_i.ifmap_regs_i._10_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ),
    .B_N(\efabless_subsystem.compute_core_i.fmap_reg_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i._01_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.ifmap_regs_i._11_  (.A(\efabless_subsystem.compute_core_i.ifmap_regs_i._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i.o_ready ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.ifmap_regs_i._14_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.ifmap_regs_i._03_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.ifmap_regs_i._15_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.ifmap_regs_i._04_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.ifmap_regs_i._16_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.ifmap_regs_i._05_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.ifmap_regs_i._17_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.ifmap_regs_i._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._07_  (.A(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._08_  (.A(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_core_i.ifmap_regs_i._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_core_i.fmap_reg_valid ),
    .A1(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_d ),
    .S(\efabless_subsystem.compute_core_i.ifmap_regs_i._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.ifmap_regs_i._05_ ),
    .S(\efabless_subsystem.compute_core_i.ifmap_regs_i._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._11_  (.A(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.fmap_reg_valid ),
    .Q_N(\efabless_subsystem.compute_core_i.ifmap_regs_i.data_valid_q_reg[0]._06_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.mux_152_27.g1._1_  (.A0(\efabless_subsystem.compute_core_i.mux_152_27.g1.data0 ),
    .A1(\efabless_subsystem.compute_core_i.mux_152_27.g1.data1 ),
    .S(\efabless_subsystem.compute_core_i.i_stat_cfg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.mux_152_27.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.mux_152_27.g1._2_  (.A(\efabless_subsystem.compute_core_i.mux_152_27.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.cdc_valid_reg[0].d ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i._158_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.acc_write_valid_reg.aclr ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_core_i.psum_accumulator_i._172_  (.A_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i._006_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._173_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i._006_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.i_acc_almost_done ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._175_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.psum_accumulator_i._008_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._177_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.psum_accumulator_i._010_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._179_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.psum_accumulator_i._012_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._184_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.psum_accumulator_i._017_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._185_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.psum_accumulator_i._018_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._186_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.psum_accumulator_i._019_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._199_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._032_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._201_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._034_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._202_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._035_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._203_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._036_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._208_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._041_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._209_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._042_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._210_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._043_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._211_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._212_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._045_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._213_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._214_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._215_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.psum_accumulator_i._216_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.psum_accumulator_i._049_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._3_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i._008_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._0_ ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._4_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.Z[1] ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._5_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i._008_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._1_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._6_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._0_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._2_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._7_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.Z[0] ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._3_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ),
    .B_N(\efabless_subsystem.compute_core_i.psum_accumulator_i._010_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._0_ ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._4_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ),
    .B_N(\efabless_subsystem.compute_core_i.psum_accumulator_i._032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._1_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._5_  (.A_N(\efabless_subsystem.compute_core_i.psum_accumulator_i._010_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._2_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._6_  (.A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._0_ ),
    .A2(\efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._1_ ),
    .B1(\efabless_subsystem.compute_core_i.psum_accumulator_i.gte_163_32._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.acc_done_q_reg.d ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._07_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.acc_write_valid_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._08_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i._034_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_d ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i._012_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i._035_ ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i._036_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._11_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .Q_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q_reg[0]._06_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1._1_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1.data0 ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1.data1 ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1._2_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_125_17.g1._1_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i._017_ ),
    .S(\efabless_subsystem.compute_controller_i.mux_acc_start_603_11.g1.z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_125_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_125_17.g1._2_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_125_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_132_31.g1._1_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i._041_ ),
    .S(\efabless_subsystem.compute_controller_i.acc_done_q_reg.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_132_31.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_132_31.g1._2_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_132_31.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_main_state_d_120_11.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1._1_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i._043_ ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.Z[1] ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1._2_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2._1_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i._042_ ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.Z[0] ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i.main_state_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2._2_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2.z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.acc_write_valid_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i._044_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g2.z ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i._018_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i._045_ ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i._046_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[0] ),
    .Q_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._07_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.acc_write_valid_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._08_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._00_ ),
    .B(\efabless_subsystem.compute_core_i.psum_accumulator_i._047_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._09_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i.mux_progress_cnt_d_120_11.g1.z ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i._019_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._10_  (.A0(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.psum_accumulator_i._048_ ),
    .S(\efabless_subsystem.compute_core_i.psum_accumulator_i._049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._11_  (.A(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._02_ ),
    .D(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.psum_accumulator_i.add_130_45.A[1] ),
    .Q_N(\efabless_subsystem.compute_core_i.psum_accumulator_i.progress_cnt_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i._07_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0].aclr ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i._08_  (.A0(\efabless_subsystem.compute_core_i.shftsgn_reg_valid ),
    .A1(\efabless_subsystem.compute_core_i.i_array_shftsgn_valid ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.shftsgn_regs_i._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i._09_  (.A(\efabless_subsystem.compute_core_i.shftsgn_regs_i._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_d ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i._10_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ),
    .B_N(\efabless_subsystem.compute_core_i.shftsgn_reg_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.shftsgn_regs_i._01_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i._11_  (.A(\efabless_subsystem.compute_core_i.shftsgn_regs_i._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.o_array_shftsgn_ready ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i._14_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.shftsgn_regs_i._03_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i._15_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.shftsgn_regs_i._04_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i._16_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.shftsgn_regs_i._05_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i._17_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.shftsgn_regs_i._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._07_  (.A(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._08_  (.A(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_core_i.shftsgn_regs_i._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_core_i.shftsgn_reg_valid ),
    .A1(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_d ),
    .S(\efabless_subsystem.compute_core_i.shftsgn_regs_i._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.shftsgn_regs_i._05_ ),
    .S(\efabless_subsystem.compute_core_i.shftsgn_regs_i._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._11_  (.A(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.shftsgn_reg_valid ),
    .Q_N(\efabless_subsystem.compute_core_i.shftsgn_regs_i.data_valid_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.weight_regs_i._07_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0].aclr ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.weight_regs_i._08_  (.A0(\efabless_subsystem.compute_core_i.weight_reg_valid ),
    .A1(\efabless_subsystem.compute_core_i.i_weight_valid ),
    .S(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.weight_regs_i._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.weight_regs_i._09_  (.A(\efabless_subsystem.compute_core_i.weight_regs_i._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_d ));
 sky130_fd_sc_hd__or2b_2 \efabless_subsystem.compute_core_i.weight_regs_i._10_  (.A(\efabless_subsystem.compute_core_i.cdc_gen.array_cdc_i.o_ready ),
    .B_N(\efabless_subsystem.compute_core_i.weight_reg_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.weight_regs_i._01_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.weight_regs_i._11_  (.A(\efabless_subsystem.compute_core_i.weight_regs_i._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.o_weight_ready ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.weight_regs_i._14_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.compute_core_i.weight_regs_i._03_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.weight_regs_i._15_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.weight_regs_i._04_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.weight_regs_i._16_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.weight_regs_i._05_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.compute_core_i.weight_regs_i._17_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.compute_core_i.weight_regs_i._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._07_  (.A(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._08_  (.A(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._00_ ),
    .B(\efabless_subsystem.compute_core_i.weight_regs_i._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._09_  (.A0(\efabless_subsystem.compute_core_i.weight_reg_valid ),
    .A1(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_d ),
    .S(\efabless_subsystem.compute_core_i.weight_regs_i._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._10_  (.A0(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.compute_core_i.weight_regs_i._05_ ),
    .S(\efabless_subsystem.compute_core_i.weight_regs_i._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._11_  (.A(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._02_ ),
    .D(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.weight_reg_valid ),
    .Q_N(\efabless_subsystem.compute_core_i.weight_regs_i.data_valid_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2633_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2634_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_auto_restart_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.config_regs_i._2635_  (.A_N(\efabless_subsystem.config_regs_i.start_q_prv ),
    .B(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g32.data0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0040_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2636_  (.A(\efabless_subsystem.config_regs_i._0040_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.i_start ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2637_  (.A(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.idle_q_reg.srd ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2638_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_start_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2640_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_mem_mode_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2641_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2642_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_soft_rst_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2643_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_global_ien_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2644_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_done_ien_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2645_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.ctl[0] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.config_regs_i._2646_  (.A(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g29.data0 ),
    .B(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0041_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2647_  (.A(\efabless_subsystem.config_regs_i._0041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2648_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2649_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2650_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_127.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2651_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2652_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_136.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2653_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2654_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_146.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2655_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2656_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_156.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2657_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2658_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_166.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2659_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2660_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_176.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2661_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2662_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_186.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2663_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2664_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_195.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2665_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2666_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_205.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2667_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2668_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_215.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2669_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2670_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_225.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2671_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2672_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_235.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2673_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2674_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_245.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2675_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2676_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_255.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2677_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2678_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_265.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2679_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2680_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_275.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2681_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2682_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_284.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2683_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2684_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_293.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2685_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2686_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_303.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2687_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2688_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_313.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2689_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2690_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_323.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2691_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2692_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_333.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2693_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2694_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_343.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2695_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2696_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_353.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2697_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2698_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_363.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2699_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2700_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_373.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2701_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2702_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_383.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2703_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2704_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_393.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2705_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2706_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_403.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2707_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2708_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_413.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2709_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2710_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_423.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2711_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424.out_0[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2712_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_358_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2744_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2745_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2746_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_624.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2747_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2748_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_632.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2749_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2750_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_640.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2751_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2752_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_648.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2753_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2754_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_656.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2755_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2756_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_664.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2757_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2758_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_672.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2759_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2760_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_680.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2761_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2762_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_688.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2763_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2764_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_696.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2765_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2766_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_704.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2767_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2768_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_712.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2769_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2808_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2809_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_873.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2810_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_879.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2811_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_885.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2812_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_891.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2813_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_897.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2814_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_903.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2815_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_909.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2816_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_915.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2817_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_921.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2818_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_927.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2819_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_933.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2820_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_939.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2840_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2841_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1061.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2842_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1067.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2843_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1073.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2844_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1079.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2845_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1085.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2846_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1091.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2847_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1097.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2848_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1103.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2872_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_21.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2873_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1249.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2874_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1255.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2875_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1261.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2876_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1267.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2877_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1273.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2878_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1279.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2879_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1285.ctl[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._2880_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1291.ctl[0] ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.config_regs_i._2969_  (.A_N(\efabless_subsystem.cfg_data_in[0] ),
    .B(\efabless_subsystem.config_regs_i.done_intr_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0000_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2970_  (.A(\efabless_subsystem.config_regs_i._0000_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.g1.data0 ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.config_regs_i._2973_  (.A_N(\efabless_subsystem.config_regs_i.soft_rst_q_prv ),
    .B(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g1.data0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0002_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2974_  (.A(\efabless_subsystem.config_regs_i._0002_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_controller_i.context_fsm_state_q_reg[0].srl ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2975_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0003_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2976_  (.A(\efabless_subsystem.config_regs_i._0003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2977_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0004_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2978_  (.A(\efabless_subsystem.config_regs_i._0004_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2979_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0005_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2980_  (.A(\efabless_subsystem.config_regs_i._0005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2981_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0006_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2982_  (.A(\efabless_subsystem.config_regs_i._0006_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2983_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0007_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2984_  (.A(\efabless_subsystem.config_regs_i._0007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2985_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0008_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2986_  (.A(\efabless_subsystem.config_regs_i._0008_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2987_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0009_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2988_  (.A(\efabless_subsystem.config_regs_i._0009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2989_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0010_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2990_  (.A(\efabless_subsystem.config_regs_i._0010_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2991_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0011_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2992_  (.A(\efabless_subsystem.config_regs_i._0011_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2993_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0012_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2994_  (.A(\efabless_subsystem.config_regs_i._0012_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2995_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0013_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2996_  (.A(\efabless_subsystem.config_regs_i._0013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2997_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0014_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._2998_  (.A(\efabless_subsystem.config_regs_i._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._2999_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0015_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3000_  (.A(\efabless_subsystem.config_regs_i._0015_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3001_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0016_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3002_  (.A(\efabless_subsystem.config_regs_i._0016_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3003_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0017_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3004_  (.A(\efabless_subsystem.config_regs_i._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3005_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0018_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3006_  (.A(\efabless_subsystem.config_regs_i._0018_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3007_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0019_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3008_  (.A(\efabless_subsystem.config_regs_i._0019_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3009_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0020_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3010_  (.A(\efabless_subsystem.config_regs_i._0020_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3011_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0021_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3012_  (.A(\efabless_subsystem.config_regs_i._0021_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3013_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0022_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3014_  (.A(\efabless_subsystem.config_regs_i._0022_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3015_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0023_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3016_  (.A(\efabless_subsystem.config_regs_i._0023_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3017_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0024_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3018_  (.A(\efabless_subsystem.config_regs_i._0024_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3019_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0025_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3020_  (.A(\efabless_subsystem.config_regs_i._0025_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3021_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0026_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3022_  (.A(\efabless_subsystem.config_regs_i._0026_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3023_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0027_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3024_  (.A(\efabless_subsystem.config_regs_i._0027_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3025_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0028_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3026_  (.A(\efabless_subsystem.config_regs_i._0028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3027_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0029_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3028_  (.A(\efabless_subsystem.config_regs_i._0029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3029_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0030_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3030_  (.A(\efabless_subsystem.config_regs_i._0030_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3031_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0031_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3032_  (.A(\efabless_subsystem.config_regs_i._0031_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3033_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0032_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3034_  (.A(\efabless_subsystem.config_regs_i._0032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3035_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[4] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0033_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3036_  (.A(\efabless_subsystem.config_regs_i._0033_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.ctl[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i._3037_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[2] ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0034_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3038_  (.A(\efabless_subsystem.config_regs_i._0034_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.ctl[1] ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.config_regs_i._3039_  (.A(\efabless_subsystem.cfg_done ),
    .B(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0035_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3040_  (.A(\efabless_subsystem.config_regs_i._0035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.idle_q_reg.srl ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.config_regs_i._3043_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q ),
    .B(\efabless_subsystem.config_regs_i.idle_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0036_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3044_  (.A(\efabless_subsystem.config_regs_i._0036_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_284_33.ctl ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.config_regs_i._3045_  (.A_N(\efabless_subsystem.config_regs_i.idle_q ),
    .B(\efabless_subsystem.config_regs_i.idle_d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0037_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3046_  (.A(\efabless_subsystem.config_regs_i._0037_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_intr_q_reg.srl ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i._3047_  (.A(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i._0038_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.config_regs_i._3048_  (.A1(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q ),
    .A2(\efabless_subsystem.config_regs_i._0038_ ),
    .B1(\efabless_subsystem.config_regs_i.start_q_prv ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i._3049_  (.A(\efabless_subsystem.config_regs_i.done_intr_q ),
    .B(\efabless_subsystem.config_regs_i.global_ien_q ),
    .C(\efabless_subsystem.config_regs_i.done_ien_q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i._0039_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i._3050_  (.A(\efabless_subsystem.config_regs_i._0039_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.o_doneintr ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i._3051_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mux_rden_198_21.ctl ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3054_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3088_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0078_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3089_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3090_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3093_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0083_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3094_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0084_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3095_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0085_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3096_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0086_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3100_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3102_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3103_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3104_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3105_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3106_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3107_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0097_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3108_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0098_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3109_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0099_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3110_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0100_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3111_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0101_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3112_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0102_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3113_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3114_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0104_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3115_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0105_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3116_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0106_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3117_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0107_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3118_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0108_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3119_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0109_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3120_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0110_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3121_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3122_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0112_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3123_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0113_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3124_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0114_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3125_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0115_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3126_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0116_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3127_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0117_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3128_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0118_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3129_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0119_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3130_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0120_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3131_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0121_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3132_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0122_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3133_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0123_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3134_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0124_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3135_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0125_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3136_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0126_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3137_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0127_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3169_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0159_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3170_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0160_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3171_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0161_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3172_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0162_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3180_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0170_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3191_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0181_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3194_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0184_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3195_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0185_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3196_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0186_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3197_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0187_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3198_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0188_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3199_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0189_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3200_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0190_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3201_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0191_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3202_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0192_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3203_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0193_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3204_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0194_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3212_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0202_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3223_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0213_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3226_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0216_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3227_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0217_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3228_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0218_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3229_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0219_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3230_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0220_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3231_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0221_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3232_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0222_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3233_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0223_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3244_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0234_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3255_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0245_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3258_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0248_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3259_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0249_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3260_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0250_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3261_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0251_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3262_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0252_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3263_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0253_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3265_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0255_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3276_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0266_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3287_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0277_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3290_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0280_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3291_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0281_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3292_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0282_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3293_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0283_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3294_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0284_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3295_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0285_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3361_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0351_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3362_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0352_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3395_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0385_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3396_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.config_regs_i._0386_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3429_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0419_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3430_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0420_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3431_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0421_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3529_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0519_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3530_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0520_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3531_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0521_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3532_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0522_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3534_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0524_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3535_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0525_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3536_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0526_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3537_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0527_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3538_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0528_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3539_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0529_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3540_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0530_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3541_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0531_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3542_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0532_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3543_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0533_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3546_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0536_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3579_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0569_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3580_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0570_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3581_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0571_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3582_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0572_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3829_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0819_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3830_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0820_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3831_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0821_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3864_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0854_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3865_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0855_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3866_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0856_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3963_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0953_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3964_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0954_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3965_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0955_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3966_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0956_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3967_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0957_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3968_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0958_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3969_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0959_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3970_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0960_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3971_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0961_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3972_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0962_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3973_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0963_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3974_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0964_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3975_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0965_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3976_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0966_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3977_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0967_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3978_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0968_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3979_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0969_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3980_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0970_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3981_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0971_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3982_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0972_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3983_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0973_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3984_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0974_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3985_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0975_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3986_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0976_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3987_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0977_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3988_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0978_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3989_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0979_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3990_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0980_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3991_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0981_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3992_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0982_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3993_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0983_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3994_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0984_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3995_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0985_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3996_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0986_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3997_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0987_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3998_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0988_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._3999_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0989_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4000_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0990_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4001_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0991_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4002_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0992_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4003_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0993_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4004_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0994_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4005_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0995_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4006_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0996_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4007_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0997_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4008_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0998_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4009_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._0999_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4010_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1000_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4011_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1001_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4012_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1002_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4013_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1003_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4014_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1004_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4015_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1005_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4016_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1006_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4017_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1007_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4018_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1008_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4019_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1009_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4020_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1010_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4021_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1011_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4022_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1012_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4023_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1013_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4024_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1014_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4025_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1015_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4026_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1016_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4027_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1017_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4028_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1018_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4029_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1019_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4030_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1020_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4031_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1021_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4032_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1022_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4033_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1023_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4034_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1024_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4035_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1025_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4036_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1026_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4037_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1027_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4038_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1028_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4039_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1029_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4040_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1030_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4041_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1031_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4042_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1032_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4043_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1033_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4044_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1034_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4045_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1035_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4046_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1036_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4047_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1037_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4048_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1038_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4049_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1039_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4050_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1040_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4051_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1041_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4052_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1042_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4053_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1043_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4054_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4055_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1045_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4056_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4057_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4058_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4059_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1049_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4060_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1050_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4061_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1051_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4062_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1052_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4063_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1053_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4064_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1054_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4065_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1055_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4066_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1056_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4067_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1057_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4068_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1058_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4069_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1059_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4070_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1060_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4071_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1061_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4072_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1062_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4073_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1063_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4074_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1064_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4075_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1065_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4076_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1066_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4077_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1067_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4078_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1068_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4079_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1069_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4080_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1070_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4081_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1071_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4082_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1072_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4083_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1073_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4084_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1074_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4085_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1075_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4086_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1076_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4087_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1077_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4088_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1078_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4089_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4090_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4091_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1081_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4092_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1082_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4093_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1083_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4094_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1084_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4095_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1085_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4096_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1086_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4097_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1087_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4098_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1088_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4099_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1089_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4100_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4101_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1091_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4102_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4103_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4104_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4105_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4106_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4107_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1097_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4108_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1098_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4109_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1099_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4110_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1100_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4111_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1101_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4112_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1102_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4113_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4114_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1104_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4115_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1105_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4116_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1106_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4117_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1107_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4118_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1108_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4119_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1109_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4120_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1110_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4121_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4122_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1112_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4123_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1113_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4124_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1114_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4125_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1115_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4126_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1116_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4127_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1117_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4128_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1118_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4129_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1119_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4130_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1120_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4131_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1121_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4132_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1122_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4133_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1123_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4134_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1124_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4135_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1125_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4136_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1126_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4137_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1127_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4138_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1128_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4139_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1129_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4140_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1130_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4141_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1131_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4142_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1132_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4143_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1133_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4144_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1134_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4145_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1135_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4146_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1136_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4147_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1137_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4148_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1138_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4149_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1139_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4150_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1140_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4151_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1141_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4152_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1142_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4153_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1143_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4154_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1144_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4155_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1145_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4156_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1146_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4157_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1147_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4158_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1148_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4159_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1149_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4160_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1150_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4161_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1151_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4255_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1245_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4256_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1246_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4257_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1247_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4258_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1248_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4259_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1249_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4260_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1250_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4261_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1251_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4262_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1252_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4263_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1253_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4264_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1254_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4265_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1255_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4266_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1256_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4288_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1278_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4289_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1279_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4290_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1280_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4321_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1311_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4322_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1312_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4323_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1313_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4330_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1320_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4331_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1321_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4332_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1322_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4333_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1323_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4334_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1324_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4335_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1325_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4336_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1326_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4337_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1327_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4338_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1328_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4339_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1329_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4340_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1330_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4341_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1331_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4342_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1332_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4343_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1333_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4344_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1334_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4345_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1335_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4346_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1336_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4347_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1337_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4348_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1338_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4349_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1339_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4350_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1340_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4351_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1341_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4352_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1342_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4353_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1343_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4354_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1344_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4355_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1345_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4356_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1346_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4357_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1347_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4358_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1348_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4359_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1349_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4360_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1350_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4361_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1351_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4362_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1352_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4384_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1374_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4385_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1375_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4386_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1376_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4417_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1407_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4418_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1408_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4419_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1409_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4426_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1416_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4427_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1417_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4428_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1418_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4429_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1419_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4430_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1420_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4431_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1421_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4432_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1422_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4433_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1423_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4434_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1424_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4435_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1425_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4436_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1426_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4437_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1427_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4438_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1428_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4439_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1429_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4440_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1430_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4441_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1431_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4442_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1432_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4443_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1433_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4444_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1434_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4445_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1435_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4446_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1436_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4447_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1437_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4448_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1438_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4449_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1439_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4480_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1470_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4481_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1471_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4482_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1472_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4513_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1503_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4514_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1504_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4515_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1505_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4522_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1512_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4523_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1513_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4524_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1514_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4525_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1515_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4526_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1516_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4527_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1517_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4528_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1518_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4529_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1519_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4530_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1520_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4531_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1521_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4532_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1522_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4533_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1523_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4534_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1524_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4535_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1525_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4536_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1526_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4537_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1527_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4538_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1528_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4539_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1529_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4543_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1533_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4544_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1534_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4545_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1535_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4576_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1566_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4577_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1567_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4578_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1568_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4609_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1599_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4610_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1600_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4611_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1601_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4618_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1608_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4619_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1609_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4620_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1610_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4621_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1611_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4622_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1612_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4623_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1613_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4624_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1614_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4625_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1615_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4626_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1616_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4627_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1617_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4628_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1618_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4629_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1619_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4630_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1620_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4631_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1621_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4632_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1622_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4633_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1623_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4634_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1624_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4635_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1625_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4831_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1821_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4832_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1822_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4833_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1823_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4834_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1824_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4835_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1825_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4836_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1826_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4837_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1827_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4838_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1828_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4839_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1829_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4840_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1830_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4841_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1831_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4842_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1832_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4864_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1854_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4865_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1855_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4866_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1856_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4897_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1887_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4898_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1888_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4899_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1889_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4906_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1896_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4907_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1897_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4908_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1898_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4909_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1899_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4910_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1900_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4911_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1901_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4912_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1902_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4913_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1903_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4914_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1904_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4915_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1905_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4916_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1906_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4917_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1907_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4918_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1908_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4919_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1909_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4920_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1910_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4921_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1911_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4922_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1912_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4923_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1913_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4924_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1914_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4925_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1915_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4926_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1916_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4927_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1917_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4928_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1918_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4929_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1919_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4930_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1920_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4931_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1921_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4932_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1922_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4933_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1923_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4934_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1924_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4935_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1925_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4936_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1926_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4937_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1927_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4938_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1928_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4960_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1950_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4961_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1951_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4962_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1952_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4993_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1983_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4994_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1984_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._4995_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1985_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5002_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1992_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5003_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1993_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5004_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1994_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5005_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1995_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5006_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1996_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5007_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1997_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5008_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1998_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5009_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._1999_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5010_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2000_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5011_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2001_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5012_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2002_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5013_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2003_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5014_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2004_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5015_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2005_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5016_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2006_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5017_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2007_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5018_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2008_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5019_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2009_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5020_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2010_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5021_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2011_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5022_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2012_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5023_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2013_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5024_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2014_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5025_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2015_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5056_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5057_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5058_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5089_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5090_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5091_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2081_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5098_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2088_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5099_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2089_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5100_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5101_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2091_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5102_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5103_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5104_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5105_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5106_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5107_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2097_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5108_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2098_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5109_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2099_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5110_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2100_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5111_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2101_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5112_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2102_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5113_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5114_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2104_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5115_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2105_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5119_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2109_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5120_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2110_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5121_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5152_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2142_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5153_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2143_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5154_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2144_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5185_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2175_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5186_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2176_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5187_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2177_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5194_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2184_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5195_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2185_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5196_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2186_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5197_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2187_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5198_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2188_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5199_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2189_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5200_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2190_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5201_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2191_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5202_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2192_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5203_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2193_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5204_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2194_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5205_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2195_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5206_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2196_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5207_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2197_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5208_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2198_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5209_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2199_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5210_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2200_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5211_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2201_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5407_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2397_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5408_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2398_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5409_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2399_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5410_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2400_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5411_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2401_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5412_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2402_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5509_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2499_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5510_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2500_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5511_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2501_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5512_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2502_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5513_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2503_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.config_regs_i._5514_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.config_regs_i._2504_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.auto_restart_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.auto_restart_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.auto_restart_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.auto_restart_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.auto_restart_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.auto_restart_q ),
    .A1(\efabless_subsystem.config_regs_i.auto_restart_d ),
    .S(\efabless_subsystem.config_regs_i._0044_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.auto_restart_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.auto_restart_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.auto_restart_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0420_ ),
    .S(\efabless_subsystem.config_regs_i._0421_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.auto_restart_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.auto_restart_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.auto_restart_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.auto_restart_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.auto_restart_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.auto_restart_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.auto_restart_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.auto_restart_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.auto_restart_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.auto_restart_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.auto_restart_q ),
    .Q_N(\efabless_subsystem.config_regs_i.auto_restart_q_reg._06_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED3 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED3 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED5 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED5 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED7 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED7 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED9 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED9 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED11 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED11 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED13 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED13 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED15 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED15 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED17 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED17 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED19 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED19 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED1 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._11_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._04_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._12_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21._04_ ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[1] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED21 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED21 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED23 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED23 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED25 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED25 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED27 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED27 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED29 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED29 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED31 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED31 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED33 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED33 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED35 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED35 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED37 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED37 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED39 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED39 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED41 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED41 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED43 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED43 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED45 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED45 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED47 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED47 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED49 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED49 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED51 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED51 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED53 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED53 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED55 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED55 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED57 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED57 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED59 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED59 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED61 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED61 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._05_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._06_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._07_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._08_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._03_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._09_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.UNCONNECTED63 ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421._10_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.UNCONNECTED63 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421.out_0[2] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[5] ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._20_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._05_ ),
    .C(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._21_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[4] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._22_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._05_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[3] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[5] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[5] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[5] ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._11_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._12_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._01_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._13_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._14_  (.A(\efabless_subsystem.cfg_address[4] ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._01_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._15_  (.A(\efabless_subsystem.cfg_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._04_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._16_  (.A(\efabless_subsystem.cfg_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._05_ ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._17_  (.A_N(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._03_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._06_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._18_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[6] ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._19_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._05_ ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[5] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._1_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._4_  (.A(\efabless_subsystem.cfg_address[16] ),
    .B(\efabless_subsystem.cfg_address[18] ),
    .C(\efabless_subsystem.cfg_address[19] ),
    .D_N(\efabless_subsystem.cfg_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._2_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[2] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._8_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26._2_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414.out_0[2] ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424._3_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D_N(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424._1_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424._7_  (.A(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424._1_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_140._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_140._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_150._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_150._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_160._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_160._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_170._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_170._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_180._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_180._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_199._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_199._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_209._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_209._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_21._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_21._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_219._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_219._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_229._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_229._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_239._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_239._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_249._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_249._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_259._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_259._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_269._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_269._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_297._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_297._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_307._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_307._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_317._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_317._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_327._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_327._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_337._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_337._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_347._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_347._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_357._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_357._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_367._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_367._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_377._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_377._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_387._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_387._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_397._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_397._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_407._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_407._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_417._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_417._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_71._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_71._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_75._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_75._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_78._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_78._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_82._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_82._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[0] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._14_  (.A(\efabless_subsystem.cfg_address[14] ),
    .B(\efabless_subsystem.cfg_address[15] ),
    .C(\efabless_subsystem.cfg_address[13] ),
    .D(\efabless_subsystem.cfg_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._15_  (.A(\efabless_subsystem.cfg_address[18] ),
    .B(\efabless_subsystem.cfg_address[19] ),
    .C(\efabless_subsystem.cfg_address[17] ),
    .D(\efabless_subsystem.cfg_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._01_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._16_  (.A(\efabless_subsystem.cfg_address[22] ),
    .B(\efabless_subsystem.cfg_address[23] ),
    .C(\efabless_subsystem.cfg_address[21] ),
    .D(\efabless_subsystem.cfg_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._02_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._17_  (.A(\efabless_subsystem.cfg_address[10] ),
    .B(\efabless_subsystem.cfg_address[11] ),
    .C(\efabless_subsystem.cfg_address[9] ),
    .D(\efabless_subsystem.cfg_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._03_ ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._18_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._01_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._02_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._19_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._05_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._20_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._06_ ));
 sky130_fd_sc_hd__and4b_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._21_  (.A_N(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._07_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._22_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._23_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._24_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[3] ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._25_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._09_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._26_  (.A(\efabless_subsystem.cfg_address[3] ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ),
    .D(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._27_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[2] ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._28_  (.A(\efabless_subsystem.cfg_address[6] ),
    .B(\efabless_subsystem.cfg_address[7] ),
    .C(\efabless_subsystem.cfg_address[5] ),
    .D(\efabless_subsystem.cfg_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._29_  (.A(\efabless_subsystem.cfg_address[2] ),
    .B(\efabless_subsystem.cfg_address[3] ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._30_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._13_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._31_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._13_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[1] ));
 sky130_fd_sc_hd__nand3_2 \efabless_subsystem.config_regs_i.ctl_i_address_312_86._32_  (.A(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._00_ ),
    .B(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._04_ ),
    .C(\efabless_subsystem.config_regs_i.ctl_i_address_312_86._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.done_ien_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.done_ien_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.done_ien_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.done_ien_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0519_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.done_ien_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.done_ien_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.done_ien_q ),
    .A1(\efabless_subsystem.config_regs_i.done_ien_d ),
    .S(\efabless_subsystem.config_regs_i._0078_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_ien_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.done_ien_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.done_ien_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0520_ ),
    .S(\efabless_subsystem.config_regs_i._0521_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_ien_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.done_ien_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.done_ien_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_ien_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.done_ien_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.done_ien_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.done_ien_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.done_ien_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.done_ien_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.done_ien_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.done_ien_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.done_ien_q ),
    .Q_N(\efabless_subsystem.config_regs_i.done_ien_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.done_intr_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.done_intr_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.done_intr_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.done_intr_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0522_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.done_intr_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.done_intr_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.done_intr_q ),
    .A1(\efabless_subsystem.config_regs_i.done_intr_d ),
    .S(\efabless_subsystem.config_regs_i._0079_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_intr_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.done_intr_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.done_intr_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0080_ ),
    .S(\efabless_subsystem.config_regs_i.done_intr_q_reg.srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_intr_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.done_intr_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.done_intr_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_intr_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.done_intr_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.done_intr_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.done_intr_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.done_intr_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.done_intr_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.done_intr_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.done_intr_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.done_intr_q ),
    .Q_N(\efabless_subsystem.config_regs_i.done_intr_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._08_  (.A(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0524_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._09_  (.A0(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv ),
    .A1(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q ),
    .S(\efabless_subsystem.config_regs_i._0083_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._10_  (.A0(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0525_ ),
    .S(\efabless_subsystem.config_regs_i._0526_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._11_  (.A(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv ),
    .Q_N(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_prv_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0527_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q ),
    .A1(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg.d ),
    .S(\efabless_subsystem.config_regs_i._0084_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0528_ ),
    .S(\efabless_subsystem.config_regs_i._0529_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q ),
    .Q_N(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.global_ien_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.global_ien_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.global_ien_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.global_ien_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0530_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.global_ien_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.global_ien_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.global_ien_q ),
    .A1(\efabless_subsystem.config_regs_i.global_ien_d ),
    .S(\efabless_subsystem.config_regs_i._0085_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.global_ien_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.global_ien_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.global_ien_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0531_ ),
    .S(\efabless_subsystem.config_regs_i._0532_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.global_ien_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.global_ien_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.global_ien_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.global_ien_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.global_ien_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.global_ien_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.global_ien_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.global_ien_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.global_ien_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.global_ien_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.global_ien_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.global_ien_q ),
    .Q_N(\efabless_subsystem.config_regs_i.global_ien_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.idle_q_reg._07_  (.A(\efabless_subsystem.config_regs_i._0533_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.idle_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.idle_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.idle_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.idle_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.idle_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.idle_q ),
    .A1(\efabless_subsystem.config_regs_i.idle_q ),
    .S(\efabless_subsystem.config_regs_i._0086_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.idle_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.idle_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.idle_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i.idle_q_reg.srd ),
    .S(\efabless_subsystem.config_regs_i.idle_q_reg.srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.idle_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.idle_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.idle_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.idle_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.idle_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.idle_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.idle_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.idle_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.idle_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.idle_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.idle_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.idle_q ),
    .Q_N(\efabless_subsystem.config_regs_i.idle_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.mem_mode_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mem_mode_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.mem_mode_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.mem_mode_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._0536_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mem_mode_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mem_mode_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .A1(\efabless_subsystem.config_regs_i.mem_mode_d ),
    .S(\efabless_subsystem.config_regs_i._0090_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mem_mode_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mem_mode_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.mem_mode_q_reg._04_ ),
    .A1(\efabless_subsystem.compute_controller_i.i_start ),
    .S(\efabless_subsystem.config_regs_i.idle_q_reg.srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mem_mode_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mem_mode_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.mem_mode_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mem_mode_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.mem_mode_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.mem_mode_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.mem_mode_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.mem_mode_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.mem_mode_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.mem_mode_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.mem_mode_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .Q_N(\efabless_subsystem.config_regs_i.mem_mode_q_reg._06_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.auto_restart_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.auto_restart_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.auto_restart_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_auto_restart_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[7] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.auto_restart_q ),
    .B2(\efabless_subsystem.config_regs_i.mux_auto_restart_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_auto_restart_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.done_ien_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_ien_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.done_ien_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_ien_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_done_ien_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.done_ien_q ),
    .B2(\efabless_subsystem.config_regs_i.mux_done_ien_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_ien_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.done_intr_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.done_intr_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.done_intr_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_intr_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.done_intr_q ),
    .B2(\efabless_subsystem.config_regs_i.mux_done_intr_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_done_intr_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i._0569_ ),
    .A1(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.fifo_ptrs_set_q_reg.d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i._0570_ ),
    .A1(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[17] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i._0571_ ),
    .B2(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_fifo_ptrs_set_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.global_ien_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.global_ien_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.global_ien_q ),
    .A1(\efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_global_ien_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_global_ien_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.global_ien_q ),
    .B2(\efabless_subsystem.config_regs_i.mux_global_ien_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_global_ien_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i._0572_ ),
    .S(\efabless_subsystem.compute_controller_i.i_start ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.idle_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_idle_d_379_18.g1._1_  (.A0(\efabless_subsystem.config_regs_i.idle_q ),
    .A1(\efabless_subsystem.config_regs_i._0092_ ),
    .S(\efabless_subsystem.cfg_done ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_idle_d_379_18.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_idle_d_379_18.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_idle_d_379_18.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_idle_d_375_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .A1(\efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mem_mode_d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .A1(\efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_mem_mode_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_mem_mode_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[16] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .B2(\efabless_subsystem.config_regs_i.mux_mem_mode_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_mem_mode_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_133.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_143.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_153.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_163.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_173.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_183.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_192.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_202.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_17.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_212.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_222.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_232.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_242.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_249.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_252.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_259.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_262.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_269.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_272.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_78.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_281.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_82.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_290.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_297.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_300.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_307.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_310.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_317.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_320.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_327.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_330.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_337.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_340.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_347.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_350.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_357.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_360.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_367.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_370.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_377.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_380.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_387.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_390.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_397.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_400.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_407.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_410.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_417.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_420.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_306_429.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_246.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_251.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_256.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_261.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_266.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_271.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_276.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_280.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_285.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_289.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_294.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_299.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_304.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_309.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_314.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_319.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_324.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_329.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_334.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_339.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_344.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_349.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_354.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_359.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_364.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_369.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_374.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_379.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_384.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_389.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_394.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_399.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_404.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_409.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_414.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_419.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_424.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_428.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_127.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[1] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_125.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_127.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_130.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_136.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[2] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_134.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_136.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_139.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_146.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[3] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_144.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_146.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_149.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_156.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[4] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_154.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_156.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_159.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_166.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[5] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_164.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_166.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_169.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_176.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[6] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_174.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_176.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_179.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_186.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[7] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_184.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_186.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_189.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_195.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[8] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_193.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_195.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_198.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_205.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[9] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_203.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_205.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_208.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_215.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[10] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_213.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_215.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_218.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_225.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[11] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_223.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_225.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_228.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_235.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[12] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_233.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_235.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_238.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_245.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[13] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_243.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_245.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_248.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_255.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[14] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_253.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_255.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_258.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_265.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[15] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_263.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_265.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_268.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_275.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[16] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_273.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_275.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_278.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_284.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[17] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_282.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_284.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_287.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_293.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[18] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_291.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_293.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_296.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_303.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[19] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_301.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_303.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_306.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_313.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[20] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_311.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_313.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_316.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_323.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[21] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_321.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_323.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_326.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_333.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[22] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_331.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_333.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_336.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_343.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[23] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_341.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_343.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_346.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_353.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[24] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_351.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_353.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_356.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_363.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[25] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_361.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_363.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_366.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_373.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[26] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_371.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_373.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_376.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_383.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[27] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_381.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_383.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_386.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_393.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[28] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_391.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_393.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_396.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_403.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[29] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_401.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_403.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_406.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_413.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[30] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_411.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_413.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_416.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_423.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[31] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_421.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_358_423.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_426.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_312_21.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_306_17.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_357_26.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_357_26.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[2] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_357_26.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_312_21.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_core_d[1]_358_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_358_21.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_358_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_357_26.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_21.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_17.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_628.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_628.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_629.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_636.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_636.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_637.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_644.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_644.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_645.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_652.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_652.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_653.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_660.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_660.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_661.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_668.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_668.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_669.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_676.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_676.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_677.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_684.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_684.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_685.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_692.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_692.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_693.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_700.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_700.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_701.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_708.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_708.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_709.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_716.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_716.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_306_717.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_21.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_628.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_636.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_644.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_652.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_660.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_668.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_676.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_684.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_692.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_700.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_708.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_312_716.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_624.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[1] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_624.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_632.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[2] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_632.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_640.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[3] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_640.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_648.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[4] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_648.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_656.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[5] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_656.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_664.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[6] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_664.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_672.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[7] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_672.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_680.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[8] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_680.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_688.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[9] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_688.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_696.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[10] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_696.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_704.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[11] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_704.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_712.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[12] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[6] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_366_712.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_21.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_17.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_876.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_876.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_877.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_882.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_882.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_883.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_888.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_888.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_889.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_894.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_894.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_895.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_900.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_900.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_901.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_906.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_906.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_907.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_912.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_912.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_913.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_918.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_918.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_919.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_924.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_211.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_924.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_209.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_925.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_930.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_221.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_930.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_219.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_931.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_936.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_231.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_936.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_229.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_937.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_942.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_241.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_942.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_239.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_306_943.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_26.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_26.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_21.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_874.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_874.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_876.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_880.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_880.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_882.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_886.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_886.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_888.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_892.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_892.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_894.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_898.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_898.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_900.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_904.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_904.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_906.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_910.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_910.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_912.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_916.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_916.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_918.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_922.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_922.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_206.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_690.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_924.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_928.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_928.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_216.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_698.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_930.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_934.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_934.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_226.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_706.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_936.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_940.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_940.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_236.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_714.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_312_942.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_26.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_873.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[1] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_873.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_874.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_879.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[2] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_879.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_880.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_885.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[3] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_885.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_886.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_891.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[4] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_891.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_892.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_897.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[5] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_897.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_898.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_903.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[6] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_903.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_904.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_909.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[7] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_909.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_910.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_915.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[8] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_915.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_916.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_921.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[9] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_686.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_921.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_922.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_927.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[10] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_694.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_927.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_928.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_933.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[11] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_702.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_933.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_934.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_939.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[12] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_710.out_0[5] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_366_939.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_357_940.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1064.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1064.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1065.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1070.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1070.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1071.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1076.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1076.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1077.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1082.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1082.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1083.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1088.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1088.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1089.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1094.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1094.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1095.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1100.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1100.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1101.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1106.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1106.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_1107.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_21.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_306_17.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1062.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1062.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1064.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1068.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1068.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1070.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1074.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1074.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1076.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1080.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1080.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1082.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1086.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1086.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1088.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1092.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1092.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1094.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1098.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1098.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1100.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1104.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1104.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_1106.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_26.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_26.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_312_21.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1061.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[1] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1061.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1062.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1067.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[2] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1067.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1068.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1073.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[3] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1073.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1074.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1079.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[4] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1079.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1080.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1085.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[5] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1085.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1086.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1091.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[6] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1091.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1092.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1097.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[7] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1097.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1098.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1103.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[8] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_1103.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_1104.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_366_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_357_26.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1252.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_132.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1252.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_75.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1253.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1258.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_142.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1258.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_140.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1259.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1264.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_152.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1264.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_150.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1265.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1270.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_162.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1270.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_160.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1271.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1276.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_172.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1276.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_170.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1277.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1282.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_182.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1282.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_180.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1283.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1288.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_191.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1288.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_21.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1289.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1294.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_201.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1294.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_199.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_1295.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_21.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .A2(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_312_21.ctl[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_21.g1.data1 ),
    .B2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_306_17.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1250.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1250.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_128.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_626.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1252.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1256.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1256.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_137.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_634.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1258.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1262.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1262.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_147.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_642.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1264.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1268.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1268.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_157.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_650.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1270.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1274.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1274.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_167.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_658.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1276.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1280.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1280.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_177.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_666.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1282.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1286.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1286.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_187.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_674.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1288.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1292.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1292.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_196.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_682.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_1294.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_26.g1._0_  (.A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_26.g1.data0 ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_offset_357_26.out_0[1] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_357_26.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_312_21.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1249.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[1] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_622.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1249.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1250.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1255.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[2] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_630.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1255.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1256.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1261.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[3] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_638.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1261.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1262.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1267.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[4] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_646.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1267.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1268.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1273.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[5] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_654.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1273.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1274.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1279.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[6] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_662.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1279.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1280.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1285.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[7] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_670.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1285.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1286.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1291.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[8] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_678.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_1291.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_1292.g1.data0 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_addressing_idx_366_21.out_0[3] ),
    .B1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .B2(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_366_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_357_26.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i._0819_ ),
    .A1(\efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i._0820_ ),
    .A1(\efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_soft_rst_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[31] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_86.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i._0821_ ),
    .B2(\efabless_subsystem.config_regs_i.mux_soft_rst_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_soft_rst_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_start_d_281_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i._0854_ ),
    .S(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g32.data0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_start_d_281_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_start_d_284_33.g1._1_  (.A0(\efabless_subsystem.config_regs_i._0855_ ),
    .A1(\efabless_subsystem.config_regs_i._0093_ ),
    .S(\efabless_subsystem.config_regs_i.mux_start_d_284_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_284_33.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_start_d_284_33.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_start_d_284_33.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_start_d_302_9.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.z ),
    .A1(\efabless_subsystem.config_regs_i.mux_start_d_302_9.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_302_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_start_d_302_9.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_start_d_302_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_302_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_start_d_306_17.g1._1_  (.A0(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.z ),
    .A1(\efabless_subsystem.config_regs_i.mux_start_d_306_17.g1.data1 ),
    .S(\efabless_subsystem.cfg_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_306_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_start_d_306_17.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_start_d_306_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_302_9.g1.data1 ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.config_regs_i.mux_start_d_312_21.g1._0_  (.A1(\efabless_subsystem.cfg_data_in[0] ),
    .A2(\efabless_subsystem.config_regs_i.ctl_i_address_312_71.out_0[4] ),
    .B1(\efabless_subsystem.config_regs_i.mux_start_d_281_9.g1.z ),
    .B2(\efabless_subsystem.config_regs_i.mux_start_d_312_21.ctl[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_start_d_306_17.g1.data1 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.mux_wren_198_21.g1._1_  (.A0(\efabless_subsystem.config_regs_i._0856_ ),
    .A1(\efabless_subsystem.cfg_wren ),
    .S(\efabless_subsystem.config_regs_i.mux_rden_198_21.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_wren_198_21.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.mux_wren_198_21.g1._2_  (.A(\efabless_subsystem.config_regs_i.mux_wren_198_21.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.mux_auto_restart_d_302_9.ctl ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ready_q_reg._07_  (.A(\efabless_subsystem.config_regs_i._0953_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ready_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.ready_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.ready_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ready_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.ready_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g29.data0 ),
    .S(\efabless_subsystem.config_regs_i._0094_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ready_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.ready_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.ready_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i.idle_q_reg.srd ),
    .S(\efabless_subsystem.config_regs_i.idle_q_reg.srl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ready_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.ready_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.ready_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.ready_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.ready_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.ready_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.ready_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.ready_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.ready_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.ready_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.ready_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g29.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.ready_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0954_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[0] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0955_ ),
    .S(\efabless_subsystem.config_regs_i._0956_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[0] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0957_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[10] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0958_ ),
    .S(\efabless_subsystem.config_regs_i._0959_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[10] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0960_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[11] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0961_ ),
    .S(\efabless_subsystem.config_regs_i._0962_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[11] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0963_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[12] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0964_ ),
    .S(\efabless_subsystem.config_regs_i._0965_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[12] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0966_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[13] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0967_ ),
    .S(\efabless_subsystem.config_regs_i._0968_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[13] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][13]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0969_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[14] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0970_ ),
    .S(\efabless_subsystem.config_regs_i._0971_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[14] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][14]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0972_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[15] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0973_ ),
    .S(\efabless_subsystem.config_regs_i._0974_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[15] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][15]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0975_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0976_ ),
    .S(\efabless_subsystem.config_regs_i._0977_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[0] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][16]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0978_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[1] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0979_ ),
    .S(\efabless_subsystem.config_regs_i._0980_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[1] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][17]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0981_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0982_ ),
    .S(\efabless_subsystem.config_regs_i._0983_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[2] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][18]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0984_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0985_ ),
    .S(\efabless_subsystem.config_regs_i._0986_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[3] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][19]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0987_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[1] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0988_ ),
    .S(\efabless_subsystem.config_regs_i._0989_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[1] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0990_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0991_ ),
    .S(\efabless_subsystem.config_regs_i._0992_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[4] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][20]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0993_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0994_ ),
    .S(\efabless_subsystem.config_regs_i._0995_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[5] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][21]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0996_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._0997_ ),
    .S(\efabless_subsystem.config_regs_i._0998_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[6] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][22]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._00_ ),
    .B(\efabless_subsystem.config_regs_i._0999_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1000_ ),
    .S(\efabless_subsystem.config_regs_i._1001_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[7] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][23]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1002_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1003_ ),
    .S(\efabless_subsystem.config_regs_i._1004_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[8] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][24]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1006_ ),
    .S(\efabless_subsystem.config_regs_i._1007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[9] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][25]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1008_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1009_ ),
    .S(\efabless_subsystem.config_regs_i._1010_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[10] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][26]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1011_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1012_ ),
    .S(\efabless_subsystem.config_regs_i._1013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[11] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][27]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1015_ ),
    .S(\efabless_subsystem.config_regs_i._1016_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[12] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][28]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1018_ ),
    .S(\efabless_subsystem.config_regs_i._1019_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[13] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][29]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1020_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[2] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1021_ ),
    .S(\efabless_subsystem.config_regs_i._1022_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[2] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1023_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1024_ ),
    .S(\efabless_subsystem.config_regs_i._1025_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[14] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][30]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1026_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._09_  (.A0(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1027_ ),
    .S(\efabless_subsystem.config_regs_i._1028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gt_269_32.A[15] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][31]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[3] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1030_ ),
    .S(\efabless_subsystem.config_regs_i._1031_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[3] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[4] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1033_ ),
    .S(\efabless_subsystem.config_regs_i._1034_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[4] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1036_ ),
    .S(\efabless_subsystem.config_regs_i._1037_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[5] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1038_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1039_ ),
    .S(\efabless_subsystem.config_regs_i._1040_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[6] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[7] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1042_ ),
    .S(\efabless_subsystem.config_regs_i._1043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[7] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1044_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[8] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1045_ ),
    .S(\efabless_subsystem.config_regs_i._1046_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[8] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1047_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._09_  (.A0(\efabless_subsystem.compute_controller_i.gte_286_30.B[9] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1048_ ),
    .S(\efabless_subsystem.config_regs_i._1049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_controller_i.gte_286_30.B[9] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[0][9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1050_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._09_  (.A0(\efabless_subsystem.compute_core_i.i_stat_cfg ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1051_ ),
    .S(\efabless_subsystem.config_regs_i._1052_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.compute_core_i.i_stat_cfg ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q2_reg[1][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1053_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.z ),
    .S(\efabless_subsystem.config_regs_i._0095_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1054_ ),
    .S(\efabless_subsystem.config_regs_i._1055_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1056_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.z ),
    .S(\efabless_subsystem.config_regs_i._0096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1057_ ),
    .S(\efabless_subsystem.config_regs_i._1058_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g22.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1059_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.z ),
    .S(\efabless_subsystem.config_regs_i._0097_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1060_ ),
    .S(\efabless_subsystem.config_regs_i._1061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g21.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.z ),
    .S(\efabless_subsystem.config_regs_i._0098_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1063_ ),
    .S(\efabless_subsystem.config_regs_i._1064_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g20.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1065_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.z ),
    .S(\efabless_subsystem.config_regs_i._0099_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1066_ ),
    .S(\efabless_subsystem.config_regs_i._1067_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g19.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][13]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1068_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.z ),
    .S(\efabless_subsystem.config_regs_i._0100_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1069_ ),
    .S(\efabless_subsystem.config_regs_i._1070_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g18.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][14]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1071_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.z ),
    .S(\efabless_subsystem.config_regs_i._0101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1072_ ),
    .S(\efabless_subsystem.config_regs_i._1073_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g17.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][15]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1074_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.z ),
    .S(\efabless_subsystem.config_regs_i._0102_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1075_ ),
    .S(\efabless_subsystem.config_regs_i._1076_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g16.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][16]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1077_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.z ),
    .S(\efabless_subsystem.config_regs_i._0103_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1078_ ),
    .S(\efabless_subsystem.config_regs_i._1079_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g15.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][17]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1080_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.z ),
    .S(\efabless_subsystem.config_regs_i._0104_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1081_ ),
    .S(\efabless_subsystem.config_regs_i._1082_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g14.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][18]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1083_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.z ),
    .S(\efabless_subsystem.config_regs_i._0105_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1084_ ),
    .S(\efabless_subsystem.config_regs_i._1085_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g13.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][19]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1086_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.z ),
    .S(\efabless_subsystem.config_regs_i._0106_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1087_ ),
    .S(\efabless_subsystem.config_regs_i._1088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g31.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1089_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.z ),
    .S(\efabless_subsystem.config_regs_i._0107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1090_ ),
    .S(\efabless_subsystem.config_regs_i._1091_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g12.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][20]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1092_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.z ),
    .S(\efabless_subsystem.config_regs_i._0108_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1093_ ),
    .S(\efabless_subsystem.config_regs_i._1094_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g11.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][21]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1095_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.z ),
    .S(\efabless_subsystem.config_regs_i._0109_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1096_ ),
    .S(\efabless_subsystem.config_regs_i._1097_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g10.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][22]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1098_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.z ),
    .S(\efabless_subsystem.config_regs_i._0110_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1099_ ),
    .S(\efabless_subsystem.config_regs_i._1100_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g9.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][23]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.z ),
    .S(\efabless_subsystem.config_regs_i._0111_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1102_ ),
    .S(\efabless_subsystem.config_regs_i._1103_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g8.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][24]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1104_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.z ),
    .S(\efabless_subsystem.config_regs_i._0112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1105_ ),
    .S(\efabless_subsystem.config_regs_i._1106_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g7.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][25]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.z ),
    .S(\efabless_subsystem.config_regs_i._0113_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1108_ ),
    .S(\efabless_subsystem.config_regs_i._1109_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g6.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][26]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1110_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.z ),
    .S(\efabless_subsystem.config_regs_i._0114_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1111_ ),
    .S(\efabless_subsystem.config_regs_i._1112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g5.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][27]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1113_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.z ),
    .S(\efabless_subsystem.config_regs_i._0115_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1114_ ),
    .S(\efabless_subsystem.config_regs_i._1115_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g4.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][28]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1116_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.z ),
    .S(\efabless_subsystem.config_regs_i._0116_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1117_ ),
    .S(\efabless_subsystem.config_regs_i._1118_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g3.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][29]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1119_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.z ),
    .S(\efabless_subsystem.config_regs_i._0117_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1120_ ),
    .S(\efabless_subsystem.config_regs_i._1121_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g30.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1122_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.z ),
    .S(\efabless_subsystem.config_regs_i._0118_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1123_ ),
    .S(\efabless_subsystem.config_regs_i._1124_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g2.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][30]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1125_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.z ),
    .S(\efabless_subsystem.config_regs_i._0119_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1126_ ),
    .S(\efabless_subsystem.config_regs_i._1127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g1.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][31]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.z ),
    .S(\efabless_subsystem.config_regs_i._0120_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1129_ ),
    .S(\efabless_subsystem.config_regs_i._1130_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g29.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1131_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.z ),
    .S(\efabless_subsystem.config_regs_i._0121_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1132_ ),
    .S(\efabless_subsystem.config_regs_i._1133_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g28.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1134_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.z ),
    .S(\efabless_subsystem.config_regs_i._0122_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1135_ ),
    .S(\efabless_subsystem.config_regs_i._1136_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g27.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1137_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.z ),
    .S(\efabless_subsystem.config_regs_i._0123_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1138_ ),
    .S(\efabless_subsystem.config_regs_i._1139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g26.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1140_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.z ),
    .S(\efabless_subsystem.config_regs_i._0124_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1141_ ),
    .S(\efabless_subsystem.config_regs_i._1142_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g25.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1143_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.z ),
    .S(\efabless_subsystem.config_regs_i._0125_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1144_ ),
    .S(\efabless_subsystem.config_regs_i._1145_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g24.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1146_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.z ),
    .S(\efabless_subsystem.config_regs_i._0126_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1147_ ),
    .S(\efabless_subsystem.config_regs_i._1148_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[0]_302_9.g23.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[0][9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1149_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.z ),
    .S(\efabless_subsystem.config_regs_i._0127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1150_ ),
    .S(\efabless_subsystem.config_regs_i._1151_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_core_d[1]_302_9.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_core_q_reg[1][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1245_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[0] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1246_ ),
    .S(\efabless_subsystem.config_regs_i._1247_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[0] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1248_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[10] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1249_ ),
    .S(\efabless_subsystem.config_regs_i._1250_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[10] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[11] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1252_ ),
    .S(\efabless_subsystem.config_regs_i._1253_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[11] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1254_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[12] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1255_ ),
    .S(\efabless_subsystem.config_regs_i._1256_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[12] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1278_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[1] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1279_ ),
    .S(\efabless_subsystem.config_regs_i._1280_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[1] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1311_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[2] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1312_ ),
    .S(\efabless_subsystem.config_regs_i._1313_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[2] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1320_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[3] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1321_ ),
    .S(\efabless_subsystem.config_regs_i._1322_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[3] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1323_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[4] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1324_ ),
    .S(\efabless_subsystem.config_regs_i._1325_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[4] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1326_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[5] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1327_ ),
    .S(\efabless_subsystem.config_regs_i._1328_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[5] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1329_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[6] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1330_ ),
    .S(\efabless_subsystem.config_regs_i._1331_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[6] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1332_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[7] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1333_ ),
    .S(\efabless_subsystem.config_regs_i._1334_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[7] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1335_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[8] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1336_ ),
    .S(\efabless_subsystem.config_regs_i._1337_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[8] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1338_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[9] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1339_ ),
    .S(\efabless_subsystem.config_regs_i._1340_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[9] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[0][9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1341_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[0] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1342_ ),
    .S(\efabless_subsystem.config_regs_i._1343_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[0] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1344_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[10] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1345_ ),
    .S(\efabless_subsystem.config_regs_i._1346_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[10] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1347_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[11] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1348_ ),
    .S(\efabless_subsystem.config_regs_i._1349_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[11] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[12] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1351_ ),
    .S(\efabless_subsystem.config_regs_i._1352_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[12] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1374_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[1] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1375_ ),
    .S(\efabless_subsystem.config_regs_i._1376_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[1] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1407_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[2] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1408_ ),
    .S(\efabless_subsystem.config_regs_i._1409_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[2] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1416_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[3] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1417_ ),
    .S(\efabless_subsystem.config_regs_i._1418_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[3] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[4] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1420_ ),
    .S(\efabless_subsystem.config_regs_i._1421_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[4] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1422_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[5] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1423_ ),
    .S(\efabless_subsystem.config_regs_i._1424_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[5] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1425_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[6] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1426_ ),
    .S(\efabless_subsystem.config_regs_i._1427_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[6] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1428_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[7] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1429_ ),
    .S(\efabless_subsystem.config_regs_i._1430_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[7] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1431_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[8] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1432_ ),
    .S(\efabless_subsystem.config_regs_i._1433_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[8] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1434_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._09_  (.A0(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[9] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1435_ ),
    .S(\efabless_subsystem.config_regs_i._1436_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[9] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[1][9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1437_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[0] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1438_ ),
    .S(\efabless_subsystem.config_regs_i._1439_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[0] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1470_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[1] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1471_ ),
    .S(\efabless_subsystem.config_regs_i._1472_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[1] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1503_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[2] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1504_ ),
    .S(\efabless_subsystem.config_regs_i._1505_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[2] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1512_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[3] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1513_ ),
    .S(\efabless_subsystem.config_regs_i._1514_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[3] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1515_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[4] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1516_ ),
    .S(\efabless_subsystem.config_regs_i._1517_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[4] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1518_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[5] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1519_ ),
    .S(\efabless_subsystem.config_regs_i._1520_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[5] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1521_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[6] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1522_ ),
    .S(\efabless_subsystem.config_regs_i._1523_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[6] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1524_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[7] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1525_ ),
    .S(\efabless_subsystem.config_regs_i._1526_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[7] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1527_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[8] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1528_ ),
    .S(\efabless_subsystem.config_regs_i._1529_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[8] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[2][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1533_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[0] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1534_ ),
    .S(\efabless_subsystem.config_regs_i._1535_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[0] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1566_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[1] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1567_ ),
    .S(\efabless_subsystem.config_regs_i._1568_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[1] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1599_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[2] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1600_ ),
    .S(\efabless_subsystem.config_regs_i._1601_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[2] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1608_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[3] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1609_ ),
    .S(\efabless_subsystem.config_regs_i._1610_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[3] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1611_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[4] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1612_ ),
    .S(\efabless_subsystem.config_regs_i._1613_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[4] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1614_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[5] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1615_ ),
    .S(\efabless_subsystem.config_regs_i._1616_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[5] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1617_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[6] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1618_ ),
    .S(\efabless_subsystem.config_regs_i._1619_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[6] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1620_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[7] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1621_ ),
    .S(\efabless_subsystem.config_regs_i._1622_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[7] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1623_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._09_  (.A0(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[8] ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .S(\efabless_subsystem.config_regs_i.count_enable_q_reg.srd ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1624_ ),
    .S(\efabless_subsystem.config_regs_i._1625_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[8] ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q2_reg[3][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1821_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.z ),
    .S(\efabless_subsystem.config_regs_i._0159_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1822_ ),
    .S(\efabless_subsystem.config_regs_i._1823_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1824_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.z ),
    .S(\efabless_subsystem.config_regs_i._0160_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1825_ ),
    .S(\efabless_subsystem.config_regs_i._1826_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g22.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1827_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.z ),
    .S(\efabless_subsystem.config_regs_i._0161_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1828_ ),
    .S(\efabless_subsystem.config_regs_i._1829_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g21.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1830_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.z ),
    .S(\efabless_subsystem.config_regs_i._0162_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1831_ ),
    .S(\efabless_subsystem.config_regs_i._1832_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g20.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1854_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.z ),
    .S(\efabless_subsystem.config_regs_i._0170_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1855_ ),
    .S(\efabless_subsystem.config_regs_i._1856_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g31.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1887_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.z ),
    .S(\efabless_subsystem.config_regs_i._0181_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1888_ ),
    .S(\efabless_subsystem.config_regs_i._1889_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g30.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1896_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.z ),
    .S(\efabless_subsystem.config_regs_i._0184_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1897_ ),
    .S(\efabless_subsystem.config_regs_i._1898_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g29.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1899_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.z ),
    .S(\efabless_subsystem.config_regs_i._0185_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1900_ ),
    .S(\efabless_subsystem.config_regs_i._1901_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g28.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1902_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.z ),
    .S(\efabless_subsystem.config_regs_i._0186_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1903_ ),
    .S(\efabless_subsystem.config_regs_i._1904_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g27.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1905_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.z ),
    .S(\efabless_subsystem.config_regs_i._0187_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1906_ ),
    .S(\efabless_subsystem.config_regs_i._1907_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g26.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1908_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.z ),
    .S(\efabless_subsystem.config_regs_i._0188_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1909_ ),
    .S(\efabless_subsystem.config_regs_i._1910_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g25.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1911_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.z ),
    .S(\efabless_subsystem.config_regs_i._0189_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1912_ ),
    .S(\efabless_subsystem.config_regs_i._1913_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g24.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1914_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.z ),
    .S(\efabless_subsystem.config_regs_i._0190_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1915_ ),
    .S(\efabless_subsystem.config_regs_i._1916_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[0]_302_9.g23.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[0][9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1917_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.z ),
    .S(\efabless_subsystem.config_regs_i._0191_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1918_ ),
    .S(\efabless_subsystem.config_regs_i._1919_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1920_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.z ),
    .S(\efabless_subsystem.config_regs_i._0192_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1921_ ),
    .S(\efabless_subsystem.config_regs_i._1922_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g22.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1923_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.z ),
    .S(\efabless_subsystem.config_regs_i._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1924_ ),
    .S(\efabless_subsystem.config_regs_i._1925_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g21.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1926_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.z ),
    .S(\efabless_subsystem.config_regs_i._0194_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1927_ ),
    .S(\efabless_subsystem.config_regs_i._1928_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g20.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1950_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.z ),
    .S(\efabless_subsystem.config_regs_i._0202_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1951_ ),
    .S(\efabless_subsystem.config_regs_i._1952_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g31.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1983_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.z ),
    .S(\efabless_subsystem.config_regs_i._0213_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1984_ ),
    .S(\efabless_subsystem.config_regs_i._1985_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g30.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1992_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.z ),
    .S(\efabless_subsystem.config_regs_i._0216_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1993_ ),
    .S(\efabless_subsystem.config_regs_i._1994_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g29.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1995_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.z ),
    .S(\efabless_subsystem.config_regs_i._0217_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1996_ ),
    .S(\efabless_subsystem.config_regs_i._1997_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g28.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._1998_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.z ),
    .S(\efabless_subsystem.config_regs_i._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._1999_ ),
    .S(\efabless_subsystem.config_regs_i._2000_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g27.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2001_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.z ),
    .S(\efabless_subsystem.config_regs_i._0219_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2002_ ),
    .S(\efabless_subsystem.config_regs_i._2003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g26.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2004_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.z ),
    .S(\efabless_subsystem.config_regs_i._0220_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2005_ ),
    .S(\efabless_subsystem.config_regs_i._2006_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g25.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.z ),
    .S(\efabless_subsystem.config_regs_i._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2008_ ),
    .S(\efabless_subsystem.config_regs_i._2009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g24.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2010_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.z ),
    .S(\efabless_subsystem.config_regs_i._0222_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2011_ ),
    .S(\efabless_subsystem.config_regs_i._2012_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[1]_302_9.g23.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[1][9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2013_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.z ),
    .S(\efabless_subsystem.config_regs_i._0223_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2014_ ),
    .S(\efabless_subsystem.config_regs_i._2015_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2046_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.z ),
    .S(\efabless_subsystem.config_regs_i._0234_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2047_ ),
    .S(\efabless_subsystem.config_regs_i._2048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g31.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2079_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.z ),
    .S(\efabless_subsystem.config_regs_i._0245_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2080_ ),
    .S(\efabless_subsystem.config_regs_i._2081_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g30.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.z ),
    .S(\efabless_subsystem.config_regs_i._0248_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2089_ ),
    .S(\efabless_subsystem.config_regs_i._2090_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g29.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2091_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.z ),
    .S(\efabless_subsystem.config_regs_i._0249_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2092_ ),
    .S(\efabless_subsystem.config_regs_i._2093_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g28.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2094_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.z ),
    .S(\efabless_subsystem.config_regs_i._0250_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2095_ ),
    .S(\efabless_subsystem.config_regs_i._2096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g27.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2097_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.z ),
    .S(\efabless_subsystem.config_regs_i._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2098_ ),
    .S(\efabless_subsystem.config_regs_i._2099_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g26.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2100_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.z ),
    .S(\efabless_subsystem.config_regs_i._0252_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2101_ ),
    .S(\efabless_subsystem.config_regs_i._2102_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g25.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2103_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.z ),
    .S(\efabless_subsystem.config_regs_i._0253_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2104_ ),
    .S(\efabless_subsystem.config_regs_i._2105_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[2]_302_9.g24.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[2][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2109_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.z ),
    .S(\efabless_subsystem.config_regs_i._0255_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2110_ ),
    .S(\efabless_subsystem.config_regs_i._2111_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2142_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.z ),
    .S(\efabless_subsystem.config_regs_i._0266_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2143_ ),
    .S(\efabless_subsystem.config_regs_i._2144_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g31.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2175_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.z ),
    .S(\efabless_subsystem.config_regs_i._0277_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2176_ ),
    .S(\efabless_subsystem.config_regs_i._2177_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g30.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2184_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.z ),
    .S(\efabless_subsystem.config_regs_i._0280_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2185_ ),
    .S(\efabless_subsystem.config_regs_i._2186_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g29.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2187_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.z ),
    .S(\efabless_subsystem.config_regs_i._0281_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2188_ ),
    .S(\efabless_subsystem.config_regs_i._2189_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g28.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2190_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.z ),
    .S(\efabless_subsystem.config_regs_i._0282_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2191_ ),
    .S(\efabless_subsystem.config_regs_i._2192_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g27.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.z ),
    .S(\efabless_subsystem.config_regs_i._0283_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2194_ ),
    .S(\efabless_subsystem.config_regs_i._2195_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g26.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2196_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.z ),
    .S(\efabless_subsystem.config_regs_i._0284_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2197_ ),
    .S(\efabless_subsystem.config_regs_i._2198_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g25.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._08_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._00_ ),
    .B(\efabless_subsystem.config_regs_i._2199_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._09_  (.A0(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.z ),
    .S(\efabless_subsystem.config_regs_i._0285_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._10_  (.A0(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2200_ ),
    .S(\efabless_subsystem.config_regs_i._2201_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._11_  (.A(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._13_  (.CLK_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._02_ ),
    .D(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_reg_mem_d[3]_302_9.g24.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.reg_mem_q_reg[3][8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._08_  (.A(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._2397_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._09_  (.A0(\efabless_subsystem.config_regs_i.soft_rst_q_prv ),
    .A1(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g1.data0 ),
    .S(\efabless_subsystem.config_regs_i._0351_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._10_  (.A0(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2398_ ),
    .S(\efabless_subsystem.config_regs_i._2399_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._11_  (.A(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.soft_rst_q_prv ),
    .Q_N(\efabless_subsystem.config_regs_i.soft_rst_q_prv_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.soft_rst_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.soft_rst_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.soft_rst_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.soft_rst_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._2400_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.soft_rst_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.soft_rst_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_soft_rst_d_302_9.g1.z ),
    .S(\efabless_subsystem.config_regs_i._0352_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.soft_rst_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.soft_rst_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.soft_rst_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2401_ ),
    .S(\efabless_subsystem.config_regs_i._2402_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.soft_rst_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.soft_rst_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.soft_rst_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.soft_rst_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.soft_rst_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.soft_rst_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.soft_rst_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.soft_rst_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.soft_rst_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.soft_rst_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.soft_rst_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g1.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.soft_rst_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.start_q_prv_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.start_q_prv_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.start_q_prv_reg._08_  (.A(\efabless_subsystem.config_regs_i.start_q_prv_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._2499_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.start_q_prv_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.start_q_prv_reg._09_  (.A0(\efabless_subsystem.config_regs_i.start_q_prv ),
    .A1(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g32.data0 ),
    .S(\efabless_subsystem.config_regs_i._0385_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.start_q_prv_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.start_q_prv_reg._10_  (.A0(\efabless_subsystem.config_regs_i.start_q_prv_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2500_ ),
    .S(\efabless_subsystem.config_regs_i._2501_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.start_q_prv_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.start_q_prv_reg._11_  (.A(\efabless_subsystem.config_regs_i.start_q_prv_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.start_q_prv_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.start_q_prv_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.start_q_prv_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.start_q_prv_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.start_q_prv_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.start_q_prv_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.start_q_prv_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.start_q_prv_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.start_q_prv ),
    .Q_N(\efabless_subsystem.config_regs_i.start_q_prv_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.start_q_reg._07_  (.A(\efabless_subsystem.config_regs_i.auto_restart_q_reg.aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.start_q_reg._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.config_regs_i.start_q_reg._08_  (.A(\efabless_subsystem.config_regs_i.start_q_reg._00_ ),
    .B(\efabless_subsystem.config_regs_i._2502_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.start_q_reg._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.start_q_reg._09_  (.A0(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g32.data0 ),
    .A1(\efabless_subsystem.config_regs_i.mux_start_d_302_9.g1.z ),
    .S(\efabless_subsystem.config_regs_i._0386_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.start_q_reg._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.config_regs_i.start_q_reg._10_  (.A0(\efabless_subsystem.config_regs_i.start_q_reg._04_ ),
    .A1(\efabless_subsystem.config_regs_i._2503_ ),
    .S(\efabless_subsystem.config_regs_i._2504_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.start_q_reg._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.config_regs_i.start_q_reg._11_  (.A(\efabless_subsystem.config_regs_i.start_q_reg._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.config_regs_i.start_q_reg._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.config_regs_i.start_q_reg._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.config_regs_i.start_q_reg._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.config_regs_i.start_q_reg._13_  (.CLK_N(\efabless_subsystem.config_regs_i.start_q_reg._02_ ),
    .D(\efabless_subsystem.config_regs_i.start_q_reg._03_ ),
    .RESET_B(\efabless_subsystem.config_regs_i.start_q_reg._00_ ),
    .SET_B(\efabless_subsystem.config_regs_i.start_q_reg._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.config_regs_i.mux_out_databuf_d_409_13.g32.data0 ),
    .Q_N(\efabless_subsystem.config_regs_i.start_q_reg._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i._162_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i._164_  (.A(\efabless_subsystem.imem_rden ),
    .B(\efabless_subsystem.input_memory_i.memory_wren ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.n_572 ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i._165_  (.A(\efabless_subsystem.input_memory_i.memory_wren ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.n_573 ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i._166_  (.A(\efabless_subsystem.imem_acc_rdata_ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i._000_ ));
 sky130_fd_sc_hd__a21o_2 \efabless_subsystem.input_memory_i._167_  (.A1(\efabless_subsystem.imem_acc_rdata_valid ),
    .A2(\efabless_subsystem.input_memory_i._000_ ),
    .B1(\efabless_subsystem.input_memory_i.eq_160_52.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.n_574 ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i._168_  (.A_N(\efabless_subsystem.input_memory_i.eq_160_52.Z ),
    .B(\efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i._001_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.input_memory_i._169_  (.A1(\efabless_subsystem.input_memory_i.eq_160_52.Z ),
    .A2(\efabless_subsystem.imem_acc_rdata_ready ),
    .A3(\efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[0] ),
    .B1(\efabless_subsystem.input_memory_i._001_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.fifo_state_reg[0].sena ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i._170_  (.A_N(\efabless_subsystem.input_memory_i.eq_159_52.Z ),
    .B(\efabless_subsystem._200_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i._002_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i._171_  (.A(\efabless_subsystem.input_memory_i._002_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_85_26.g1.data1 ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i._172_  (.A(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .B(\efabless_subsystem.input_memory_i.mux_85_26.g1.data1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i._003_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i._173_  (.A(\efabless_subsystem.input_memory_i._003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.input_memory_i._174_  (.A1(\efabless_subsystem.imem_acc_rdata_valid ),
    .A2(\efabless_subsystem.input_memory_i._000_ ),
    .B1(\efabless_subsystem.input_memory_i.eq_160_52.Z ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._175_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._010_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._176_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._011_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._177_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._012_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._178_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._013_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._179_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._014_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._180_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._015_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._181_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._016_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._182_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._017_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._183_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._018_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._184_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._019_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._185_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._020_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._186_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._021_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._187_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._022_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._188_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._023_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._189_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._024_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._190_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._025_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._191_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._026_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._192_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._027_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._193_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._028_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._194_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._029_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._195_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._030_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._196_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._031_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._197_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._032_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._198_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._033_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._199_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._034_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._200_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._035_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._201_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._036_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._202_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._037_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._203_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._038_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._204_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._039_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._205_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._040_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._206_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._041_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._207_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._042_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._208_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._043_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._209_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._210_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._045_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._211_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._212_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._213_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._214_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._049_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._215_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._050_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._216_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._051_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._217_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._052_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._218_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._053_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._219_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._054_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._220_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._055_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._221_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._056_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._222_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._057_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._223_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._058_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._224_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._059_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._225_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._060_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._226_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._061_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._227_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._062_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._228_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._063_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._229_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.input_memory_i._064_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._230_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._065_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._231_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._066_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._232_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._067_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._233_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._068_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._234_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._069_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._235_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._070_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._236_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._071_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._237_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._072_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._238_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._073_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._239_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._074_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._240_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._075_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._241_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._076_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._242_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._077_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._243_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._078_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._244_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._245_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._246_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._081_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._247_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._082_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._248_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._083_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._249_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._084_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._250_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._085_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._251_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._086_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._252_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._087_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._253_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._088_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._254_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._089_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._255_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._256_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._091_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._257_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._258_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._259_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._260_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._261_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._262_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._097_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._263_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._098_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._264_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._099_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._265_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._100_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._266_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._101_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._267_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._102_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._268_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._269_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._104_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._270_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._105_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._271_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._106_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._272_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._107_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._273_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._108_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._274_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._109_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._275_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._110_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._276_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._277_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._112_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._278_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._113_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._279_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._114_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._280_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._115_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._281_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._116_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._282_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._117_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._283_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._118_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._284_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._119_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._285_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._120_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._286_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._121_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._287_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._122_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._288_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._123_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._289_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._124_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._290_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._125_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._291_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._126_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._292_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._127_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._293_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._128_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._294_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._129_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._295_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._130_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._296_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._131_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._297_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._132_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._298_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._133_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._299_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._134_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._300_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._135_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._301_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._136_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._302_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._137_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._303_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._138_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._304_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._139_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._305_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._140_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._306_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._141_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._307_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._142_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._308_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._143_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._309_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._144_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._310_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._145_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._311_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._146_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._312_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._147_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._313_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._148_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._314_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._149_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._315_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._150_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._316_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._151_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._317_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._152_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._318_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._153_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._319_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._154_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._320_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._155_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._321_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._156_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._322_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._157_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._323_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._158_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._324_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._159_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._325_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._160_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.input_memory_i._326_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.input_memory_i._161_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_144_39._25_  (.A(\efabless_subsystem.input_memory_i._010_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .C(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_144_39._26_  (.A(\efabless_subsystem.input_memory_i.add_144_39._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._01_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.input_memory_i.add_144_39._27_  (.A1(\efabless_subsystem.input_memory_i._010_ ),
    .A2(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i.add_144_39._28_  (.A(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39.Z[1] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_144_39._29_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i.add_144_39._30_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39._04_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i.add_144_39._31_  (.A(\efabless_subsystem.input_memory_i.add_144_39._03_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39.Z[2] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_144_39._32_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_144_39._33_  (.A(\efabless_subsystem.input_memory_i.add_144_39._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._06_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.add_144_39._34_  (.A(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39._07_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.input_memory_i.add_144_39._35_  (.A1(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .A2(\efabless_subsystem.input_memory_i.add_144_39._03_ ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.input_memory_i.add_144_39._36_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39.Z[4] ));
 sky130_fd_sc_hd__nand4_2 \efabless_subsystem.input_memory_i.add_144_39._37_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .C(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .D(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39._08_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.input_memory_i.add_144_39._38_  (.A1(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .A2(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .A3(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._09_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_144_39._39_  (.A(\efabless_subsystem.input_memory_i.add_144_39._08_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_144_39._40_  (.A(\efabless_subsystem.input_memory_i.add_144_39._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[5] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.input_memory_i.add_144_39._41_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_144_39.Z[6] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_144_39._42_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .C(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .D(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_144_39._43_  (.A(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .C(\efabless_subsystem.input_memory_i.add_144_39._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_144_39._44_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .C(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._13_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.input_memory_i.add_144_39._45_  (.A1(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .A2(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .A3(\efabless_subsystem.input_memory_i.add_144_39._13_ ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._14_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i.add_144_39._46_  (.A_N(\efabless_subsystem.input_memory_i.add_144_39._12_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._15_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_144_39._47_  (.A(\efabless_subsystem.input_memory_i.add_144_39._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.add_144_39._48_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[8] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_144_39._49_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._16_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_144_39._50_  (.A(\efabless_subsystem.input_memory_i.add_144_39._00_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .C(\efabless_subsystem.input_memory_i.add_144_39._11_ ),
    .D(\efabless_subsystem.input_memory_i.add_144_39._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._17_ ));
 sky130_fd_sc_hd__a41o_2 \efabless_subsystem.input_memory_i.add_144_39._51_  (.A1(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .A2(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .A3(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .A4(\efabless_subsystem.input_memory_i.add_144_39._11_ ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._18_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i.add_144_39._52_  (.A_N(\efabless_subsystem.input_memory_i.add_144_39._17_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._19_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_144_39._53_  (.A(\efabless_subsystem.input_memory_i.add_144_39._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[9] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_144_39._54_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .C(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._20_ ));
 sky130_fd_sc_hd__o2bb2a_2 \efabless_subsystem.input_memory_i.add_144_39._55_  (.A1_N(\efabless_subsystem.input_memory_i.add_144_39._12_ ),
    .A2_N(\efabless_subsystem.input_memory_i.add_144_39._20_ ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39._17_ ),
    .B2(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[10] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_144_39._56_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .C(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .D(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._21_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_144_39._57_  (.A(\efabless_subsystem.input_memory_i.add_144_39._00_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .C(\efabless_subsystem.input_memory_i.add_144_39._11_ ),
    .D(\efabless_subsystem.input_memory_i.add_144_39._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._22_ ));
 sky130_fd_sc_hd__a41o_2 \efabless_subsystem.input_memory_i.add_144_39._58_  (.A1(\efabless_subsystem.input_memory_i.add_144_39._01_ ),
    .A2(\efabless_subsystem.input_memory_i.add_144_39._06_ ),
    .A3(\efabless_subsystem.input_memory_i.add_144_39._11_ ),
    .A4(\efabless_subsystem.input_memory_i.add_144_39._20_ ),
    .B1(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._23_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i.add_144_39._59_  (.A_N(\efabless_subsystem.input_memory_i.add_144_39._22_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._23_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39._24_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_144_39._60_  (.A(\efabless_subsystem.input_memory_i.add_144_39._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[11] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.add_144_39._61_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[12] ),
    .B(\efabless_subsystem.input_memory_i.add_144_39._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[12] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.add_144_39._62_  (.A(\efabless_subsystem.input_memory_i._010_ ),
    .B(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_144_39.Z[0] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_149_37._25_  (.A(\efabless_subsystem.input_memory_i._011_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .C(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._00_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_149_37._26_  (.A(\efabless_subsystem.input_memory_i.add_149_37._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._01_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.input_memory_i.add_149_37._27_  (.A1(\efabless_subsystem.input_memory_i._011_ ),
    .A2(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i.add_149_37._28_  (.A(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._02_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37.Z[1] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_149_37._29_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i.add_149_37._30_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37._04_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.input_memory_i.add_149_37._31_  (.A(\efabless_subsystem.input_memory_i.add_149_37._03_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37.Z[2] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_149_37._32_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_149_37._33_  (.A(\efabless_subsystem.input_memory_i.add_149_37._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._06_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.add_149_37._34_  (.A(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37._07_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.input_memory_i.add_149_37._35_  (.A1(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .A2(\efabless_subsystem.input_memory_i.add_149_37._03_ ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.input_memory_i.add_149_37._36_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37.Z[4] ));
 sky130_fd_sc_hd__nand4_2 \efabless_subsystem.input_memory_i.add_149_37._37_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .C(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .D(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37._08_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.input_memory_i.add_149_37._38_  (.A1(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .A2(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .A3(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._09_ ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_149_37._39_  (.A(\efabless_subsystem.input_memory_i.add_149_37._08_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._10_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_149_37._40_  (.A(\efabless_subsystem.input_memory_i.add_149_37._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[5] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.input_memory_i.add_149_37._41_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.add_149_37.Z[6] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_149_37._42_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .C(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .D(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._11_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_149_37._43_  (.A(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .C(\efabless_subsystem.input_memory_i.add_149_37._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._12_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_149_37._44_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .C(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._13_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.input_memory_i.add_149_37._45_  (.A1(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .A2(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .A3(\efabless_subsystem.input_memory_i.add_149_37._13_ ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._14_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i.add_149_37._46_  (.A_N(\efabless_subsystem.input_memory_i.add_149_37._12_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._14_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._15_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_149_37._47_  (.A(\efabless_subsystem.input_memory_i.add_149_37._15_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.add_149_37._48_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[8] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.input_memory_i.add_149_37._49_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._16_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_149_37._50_  (.A(\efabless_subsystem.input_memory_i.add_149_37._00_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .C(\efabless_subsystem.input_memory_i.add_149_37._11_ ),
    .D(\efabless_subsystem.input_memory_i.add_149_37._16_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._17_ ));
 sky130_fd_sc_hd__a41o_2 \efabless_subsystem.input_memory_i.add_149_37._51_  (.A1(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .A2(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .A3(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .A4(\efabless_subsystem.input_memory_i.add_149_37._11_ ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._18_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i.add_149_37._52_  (.A_N(\efabless_subsystem.input_memory_i.add_149_37._17_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._19_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_149_37._53_  (.A(\efabless_subsystem.input_memory_i.add_149_37._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[9] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.input_memory_i.add_149_37._54_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .C(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._20_ ));
 sky130_fd_sc_hd__o2bb2a_2 \efabless_subsystem.input_memory_i.add_149_37._55_  (.A1_N(\efabless_subsystem.input_memory_i.add_149_37._12_ ),
    .A2_N(\efabless_subsystem.input_memory_i.add_149_37._20_ ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37._17_ ),
    .B2(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[10] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_149_37._56_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .C(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .D(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._21_ ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.input_memory_i.add_149_37._57_  (.A(\efabless_subsystem.input_memory_i.add_149_37._00_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .C(\efabless_subsystem.input_memory_i.add_149_37._11_ ),
    .D(\efabless_subsystem.input_memory_i.add_149_37._21_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._22_ ));
 sky130_fd_sc_hd__a41o_2 \efabless_subsystem.input_memory_i.add_149_37._58_  (.A1(\efabless_subsystem.input_memory_i.add_149_37._01_ ),
    .A2(\efabless_subsystem.input_memory_i.add_149_37._06_ ),
    .A3(\efabless_subsystem.input_memory_i.add_149_37._11_ ),
    .A4(\efabless_subsystem.input_memory_i.add_149_37._20_ ),
    .B1(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._23_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.input_memory_i.add_149_37._59_  (.A_N(\efabless_subsystem.input_memory_i.add_149_37._22_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._23_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37._24_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.add_149_37._60_  (.A(\efabless_subsystem.input_memory_i.add_149_37._24_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[11] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.add_149_37._61_  (.A(\efabless_subsystem.input_memory_i.add_149_37.A[12] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37._22_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[12] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.add_149_37._62_  (.A(\efabless_subsystem.input_memory_i._011_ ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.add_149_37.Z[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.ctl_fifo_state_103_19._0_  (.A(\efabless_subsystem.imem_acc_rdata_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.input_memory_i.ctl_fifo_state_103_19._1_  (.A(\efabless_subsystem.imem_acc_rdata_valid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[0] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._20_  (.A(\efabless_subsystem.input_memory_i._065_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._00_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._21_  (.A(\efabless_subsystem.input_memory_i._069_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._01_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.eq_159_52._22_  (.A(\efabless_subsystem.input_memory_i.eq_159_52.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.eq_159_52._02_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.eq_159_52._23_  (.A(\efabless_subsystem.input_memory_i._070_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.eq_159_52._03_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._24_  (.A(\efabless_subsystem.input_memory_i._074_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._04_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.input_memory_i.eq_159_52._25_  (.A1(\efabless_subsystem.input_memory_i._012_ ),
    .A2(\efabless_subsystem.input_memory_i.eq_159_52._02_ ),
    .B1(\efabless_subsystem.input_memory_i.eq_159_52._03_ ),
    .B2(\efabless_subsystem.input_memory_i.eq_159_52.A[5] ),
    .C1(\efabless_subsystem.input_memory_i.eq_159_52._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._05_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.eq_159_52._26_  (.A(\efabless_subsystem.input_memory_i._067_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.eq_159_52._06_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.input_memory_i.eq_159_52._27_  (.A(\efabless_subsystem.input_memory_i._067_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._07_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.eq_159_52._28_  (.A(\efabless_subsystem.input_memory_i._066_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.eq_159_52._08_ ));
 sky130_fd_sc_hd__or2_2 \efabless_subsystem.input_memory_i.eq_159_52._29_  (.A(\efabless_subsystem.input_memory_i._066_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._09_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._30_  (.A(\efabless_subsystem.input_memory_i._075_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._10_ ));
 sky130_fd_sc_hd__a221o_2 \efabless_subsystem.input_memory_i.eq_159_52._31_  (.A1(\efabless_subsystem.input_memory_i.eq_159_52._06_ ),
    .A2(\efabless_subsystem.input_memory_i.eq_159_52._07_ ),
    .B1(\efabless_subsystem.input_memory_i.eq_159_52._08_ ),
    .B2(\efabless_subsystem.input_memory_i.eq_159_52._09_ ),
    .C1(\efabless_subsystem.input_memory_i.eq_159_52._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._11_ ));
 sky130_fd_sc_hd__o22a_2 \efabless_subsystem.input_memory_i.eq_159_52._32_  (.A1(\efabless_subsystem.input_memory_i._012_ ),
    .A2(\efabless_subsystem.input_memory_i.eq_159_52._02_ ),
    .B1(\efabless_subsystem.input_memory_i.eq_159_52._03_ ),
    .B2(\efabless_subsystem.input_memory_i.eq_159_52.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._12_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.input_memory_i.eq_159_52._33_  (.A(\efabless_subsystem.input_memory_i.eq_159_52._01_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52._05_ ),
    .C(\efabless_subsystem.input_memory_i.eq_159_52._11_ ),
    .D_N(\efabless_subsystem.input_memory_i.eq_159_52._12_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._13_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._34_  (.A(\efabless_subsystem.input_memory_i._068_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._14_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._35_  (.A(\efabless_subsystem.input_memory_i._071_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._15_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._36_  (.A(\efabless_subsystem.input_memory_i._072_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._16_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._37_  (.A(\efabless_subsystem.input_memory_i._076_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._17_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_159_52._38_  (.A(\efabless_subsystem.input_memory_i._073_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._18_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.input_memory_i.eq_159_52._39_  (.A(\efabless_subsystem.input_memory_i.eq_159_52._15_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52._16_ ),
    .C(\efabless_subsystem.input_memory_i.eq_159_52._17_ ),
    .D(\efabless_subsystem.input_memory_i.eq_159_52._18_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52._19_ ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.input_memory_i.eq_159_52._40_  (.A(\efabless_subsystem.input_memory_i.eq_159_52._00_ ),
    .B(\efabless_subsystem.input_memory_i.eq_159_52._13_ ),
    .C(\efabless_subsystem.input_memory_i.eq_159_52._14_ ),
    .D(\efabless_subsystem.input_memory_i.eq_159_52._19_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.eq_159_52.Z ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.eq_160_52._4_  (.A(\efabless_subsystem.input_memory_i._077_ ),
    .B(\efabless_subsystem.input_memory_i.eq_160_52.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52._0_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.input_memory_i.eq_160_52._5_  (.A(\efabless_subsystem.input_memory_i.eq_160_52.A[11] ),
    .B(\efabless_subsystem.input_memory_i.eq_160_52.A[12] ),
    .C(\efabless_subsystem.input_memory_i.eq_160_52.A[10] ),
    .D(\efabless_subsystem.input_memory_i.eq_160_52.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52._1_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.input_memory_i.eq_160_52._6_  (.A(\efabless_subsystem.input_memory_i.eq_160_52.A[3] ),
    .B(\efabless_subsystem.input_memory_i.eq_160_52.A[4] ),
    .C(\efabless_subsystem.input_memory_i.eq_160_52.A[2] ),
    .D(\efabless_subsystem.input_memory_i.eq_160_52.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52._2_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.input_memory_i.eq_160_52._7_  (.A(\efabless_subsystem.input_memory_i.eq_160_52.A[7] ),
    .B(\efabless_subsystem.input_memory_i.eq_160_52.A[8] ),
    .C(\efabless_subsystem.input_memory_i.eq_160_52.A[6] ),
    .D(\efabless_subsystem.input_memory_i.eq_160_52.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52._3_ ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.input_memory_i.eq_160_52._8_  (.A(\efabless_subsystem.input_memory_i.eq_160_52._0_ ),
    .B(\efabless_subsystem.input_memory_i.eq_160_52._1_ ),
    .C(\efabless_subsystem.input_memory_i.eq_160_52._2_ ),
    .D(\efabless_subsystem.input_memory_i.eq_160_52._3_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.eq_160_52.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._08_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._00_ ),
    .B(\efabless_subsystem.input_memory_i._078_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._09_  (.A0(\efabless_subsystem.imem_acc_rdata_valid ),
    .A1(\efabless_subsystem.input_memory_i.fifo_state_reg[0].d ),
    .S(\efabless_subsystem.input_memory_i.fifo_state_reg[0].sena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._10_  (.A0(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._079_ ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._11_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.fifo_state_reg[0]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._02_ ),
    .D(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.imem_acc_rdata_valid ),
    .Q_N(\efabless_subsystem.input_memory_i.fifo_state_reg[0]._06_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._00_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[0] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._01_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[1] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._02_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[2] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._03_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._04_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[4] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._05_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._06_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[6] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._07_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._08_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[8] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._09_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[9] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._10_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[10] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._11_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[11] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g17._12_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[12] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_159_52.A[12] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._00_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[0] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._01_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[1] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._02_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[2] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._03_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._04_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[4] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._05_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._06_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[6] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._07_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._08_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[8] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._09_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[9] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._10_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[10] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._11_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[11] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.input_memory_i.g18._12_  (.A(\efabless_subsystem.input_memory_i.add_144_39.A[12] ),
    .B(\efabless_subsystem.input_memory_i.add_149_37.A[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.eq_160_52.A[12] ));
 sky130_sram_1kbytes_1rw1r_200x48_8 \efabless_subsystem.input_memory_i.mem200  (.csb0(\efabless_subsystem.input_memory_i.n_572 ),
    .csb1(\efabless_subsystem.input_memory_i.n_574 ),
    .web0(\efabless_subsystem.input_memory_i.n_573 ),
    .clk0(wb_clk_i),
    .clk1(wb_clk_i),
    .addr0({\efabless_subsystem.input_memory_i.memory_addr[5] ,
    \efabless_subsystem.input_memory_i.memory_addr[4] ,
    \efabless_subsystem.input_memory_i.memory_addr[3] ,
    \efabless_subsystem.input_memory_i.memory_addr[2] ,
    \efabless_subsystem.input_memory_i.memory_addr[1] ,
    \efabless_subsystem.input_memory_i.memory_addr[0] }),
    .addr1({\efabless_subsystem.input_memory_i.add_149_37.A[5] ,
    \efabless_subsystem.input_memory_i.add_149_37.A[4] ,
    \efabless_subsystem.input_memory_i.add_149_37.A[3] ,
    \efabless_subsystem.input_memory_i.add_149_37.A[2] ,
    \efabless_subsystem.input_memory_i.add_149_37.A[1] ,
    \efabless_subsystem.input_memory_i.add_149_37.A[0] }),
    .din0({\efabless_subsystem.input_memory_i._082_ ,
    \efabless_subsystem.input_memory_i._081_ ,
    \efabless_subsystem.input_memory_i._080_ ,
    \efabless_subsystem.input_memory_i.memory_wdata[196] ,
    \efabless_subsystem.input_memory_i.memory_wdata[195] ,
    \efabless_subsystem.input_memory_i.memory_wdata[194] ,
    \efabless_subsystem.input_memory_i.memory_wdata[193] ,
    \efabless_subsystem.input_memory_i.memory_wdata[192] ,
    \efabless_subsystem.input_memory_i.memory_wdata[191] ,
    \efabless_subsystem.input_memory_i.memory_wdata[190] ,
    \efabless_subsystem.input_memory_i.memory_wdata[189] ,
    \efabless_subsystem.input_memory_i.memory_wdata[188] ,
    \efabless_subsystem.input_memory_i.memory_wdata[187] ,
    \efabless_subsystem.input_memory_i.memory_wdata[186] ,
    \efabless_subsystem.input_memory_i.memory_wdata[185] ,
    \efabless_subsystem.input_memory_i.memory_wdata[184] ,
    \efabless_subsystem.input_memory_i.memory_wdata[183] ,
    \efabless_subsystem.input_memory_i.memory_wdata[182] ,
    \efabless_subsystem.input_memory_i.memory_wdata[181] ,
    \efabless_subsystem.input_memory_i.memory_wdata[180] ,
    \efabless_subsystem.input_memory_i.memory_wdata[179] ,
    \efabless_subsystem.input_memory_i.memory_wdata[178] ,
    \efabless_subsystem.input_memory_i.memory_wdata[177] ,
    \efabless_subsystem.input_memory_i.memory_wdata[176] ,
    \efabless_subsystem.input_memory_i.memory_wdata[175] ,
    \efabless_subsystem.input_memory_i.memory_wdata[174] ,
    \efabless_subsystem.input_memory_i.memory_wdata[173] ,
    \efabless_subsystem.input_memory_i.memory_wdata[172] ,
    \efabless_subsystem.input_memory_i.memory_wdata[171] ,
    \efabless_subsystem.input_memory_i.memory_wdata[170] ,
    \efabless_subsystem.input_memory_i.memory_wdata[169] ,
    \efabless_subsystem.input_memory_i.memory_wdata[168] ,
    \efabless_subsystem.input_memory_i.memory_wdata[167] ,
    \efabless_subsystem.input_memory_i.memory_wdata[166] ,
    \efabless_subsystem.input_memory_i.memory_wdata[165] ,
    \efabless_subsystem.input_memory_i.memory_wdata[164] ,
    \efabless_subsystem.input_memory_i.memory_wdata[163] ,
    \efabless_subsystem.input_memory_i.memory_wdata[162] ,
    \efabless_subsystem.input_memory_i.memory_wdata[161] ,
    \efabless_subsystem.input_memory_i.memory_wdata[160] ,
    \efabless_subsystem.input_memory_i.memory_wdata[159] ,
    \efabless_subsystem.input_memory_i.memory_wdata[158] ,
    \efabless_subsystem.input_memory_i.memory_wdata[157] ,
    \efabless_subsystem.input_memory_i.memory_wdata[156] ,
    \efabless_subsystem.input_memory_i.memory_wdata[155] ,
    \efabless_subsystem.input_memory_i.memory_wdata[154] ,
    \efabless_subsystem.input_memory_i.memory_wdata[153] ,
    \efabless_subsystem.input_memory_i.memory_wdata[152] ,
    \efabless_subsystem.input_memory_i.memory_wdata[151] ,
    \efabless_subsystem.input_memory_i.memory_wdata[150] ,
    \efabless_subsystem.input_memory_i.memory_wdata[149] ,
    \efabless_subsystem.input_memory_i.memory_wdata[148] ,
    \efabless_subsystem.input_memory_i.memory_wdata[147] ,
    \efabless_subsystem.input_memory_i.memory_wdata[146] ,
    \efabless_subsystem.input_memory_i.memory_wdata[145] ,
    \efabless_subsystem.input_memory_i.memory_wdata[144] ,
    \efabless_subsystem.input_memory_i.memory_wdata[143] ,
    \efabless_subsystem.input_memory_i.memory_wdata[142] ,
    \efabless_subsystem.input_memory_i.memory_wdata[141] ,
    \efabless_subsystem.input_memory_i.memory_wdata[140] ,
    \efabless_subsystem.input_memory_i.memory_wdata[139] ,
    \efabless_subsystem.input_memory_i.memory_wdata[138] ,
    \efabless_subsystem.input_memory_i.memory_wdata[137] ,
    \efabless_subsystem.input_memory_i.memory_wdata[136] ,
    \efabless_subsystem.input_memory_i.memory_wdata[135] ,
    \efabless_subsystem.input_memory_i.memory_wdata[134] ,
    \efabless_subsystem.input_memory_i.memory_wdata[133] ,
    \efabless_subsystem.input_memory_i.memory_wdata[132] ,
    \efabless_subsystem.input_memory_i.memory_wdata[131] ,
    \efabless_subsystem.input_memory_i.memory_wdata[130] ,
    \efabless_subsystem.input_memory_i.memory_wdata[129] ,
    \efabless_subsystem.input_memory_i.memory_wdata[128] ,
    \efabless_subsystem.input_memory_i.memory_wdata[127] ,
    \efabless_subsystem.input_memory_i.memory_wdata[126] ,
    \efabless_subsystem.input_memory_i.memory_wdata[125] ,
    \efabless_subsystem.input_memory_i.memory_wdata[124] ,
    \efabless_subsystem.input_memory_i.memory_wdata[123] ,
    \efabless_subsystem.input_memory_i.memory_wdata[122] ,
    \efabless_subsystem.input_memory_i.memory_wdata[121] ,
    \efabless_subsystem.input_memory_i.memory_wdata[120] ,
    \efabless_subsystem.input_memory_i.memory_wdata[119] ,
    \efabless_subsystem.input_memory_i.memory_wdata[118] ,
    \efabless_subsystem.input_memory_i.memory_wdata[117] ,
    \efabless_subsystem.input_memory_i.memory_wdata[116] ,
    \efabless_subsystem.input_memory_i.memory_wdata[115] ,
    \efabless_subsystem.input_memory_i.memory_wdata[114] ,
    \efabless_subsystem.input_memory_i.memory_wdata[113] ,
    \efabless_subsystem.input_memory_i.memory_wdata[112] ,
    \efabless_subsystem.input_memory_i.memory_wdata[111] ,
    \efabless_subsystem.input_memory_i.memory_wdata[110] ,
    \efabless_subsystem.input_memory_i.memory_wdata[109] ,
    \efabless_subsystem.input_memory_i.memory_wdata[108] ,
    \efabless_subsystem.input_memory_i.memory_wdata[107] ,
    \efabless_subsystem.input_memory_i.memory_wdata[106] ,
    \efabless_subsystem.input_memory_i.memory_wdata[105] ,
    \efabless_subsystem.input_memory_i.memory_wdata[104] ,
    \efabless_subsystem.input_memory_i.memory_wdata[103] ,
    \efabless_subsystem.input_memory_i.memory_wdata[102] ,
    \efabless_subsystem.input_memory_i.memory_wdata[101] ,
    \efabless_subsystem.input_memory_i.memory_wdata[100] ,
    \efabless_subsystem.input_memory_i.memory_wdata[99] ,
    \efabless_subsystem.input_memory_i.memory_wdata[98] ,
    \efabless_subsystem.input_memory_i.memory_wdata[97] ,
    \efabless_subsystem.input_memory_i.memory_wdata[96] ,
    \efabless_subsystem.input_memory_i.memory_wdata[95] ,
    \efabless_subsystem.input_memory_i.memory_wdata[94] ,
    \efabless_subsystem.input_memory_i.memory_wdata[93] ,
    \efabless_subsystem.input_memory_i.memory_wdata[92] ,
    \efabless_subsystem.input_memory_i.memory_wdata[91] ,
    \efabless_subsystem.input_memory_i.memory_wdata[90] ,
    \efabless_subsystem.input_memory_i.memory_wdata[89] ,
    \efabless_subsystem.input_memory_i.memory_wdata[88] ,
    \efabless_subsystem.input_memory_i.memory_wdata[87] ,
    \efabless_subsystem.input_memory_i.memory_wdata[86] ,
    \efabless_subsystem.input_memory_i.memory_wdata[85] ,
    \efabless_subsystem.input_memory_i.memory_wdata[84] ,
    \efabless_subsystem.input_memory_i.memory_wdata[83] ,
    \efabless_subsystem.input_memory_i.memory_wdata[82] ,
    \efabless_subsystem.input_memory_i.memory_wdata[81] ,
    \efabless_subsystem.input_memory_i.memory_wdata[80] ,
    \efabless_subsystem.input_memory_i.memory_wdata[79] ,
    \efabless_subsystem.input_memory_i.memory_wdata[78] ,
    \efabless_subsystem.input_memory_i.memory_wdata[77] ,
    \efabless_subsystem.input_memory_i.memory_wdata[76] ,
    \efabless_subsystem.input_memory_i.memory_wdata[75] ,
    \efabless_subsystem.input_memory_i.memory_wdata[74] ,
    \efabless_subsystem.input_memory_i.memory_wdata[73] ,
    \efabless_subsystem.input_memory_i.memory_wdata[72] ,
    \efabless_subsystem.input_memory_i.memory_wdata[71] ,
    \efabless_subsystem.input_memory_i.memory_wdata[70] ,
    \efabless_subsystem.input_memory_i.memory_wdata[69] ,
    \efabless_subsystem.input_memory_i.memory_wdata[68] ,
    \efabless_subsystem.input_memory_i.memory_wdata[67] ,
    \efabless_subsystem.input_memory_i.memory_wdata[66] ,
    \efabless_subsystem.input_memory_i.memory_wdata[65] ,
    \efabless_subsystem.input_memory_i.memory_wdata[64] ,
    \efabless_subsystem.input_memory_i.memory_wdata[63] ,
    \efabless_subsystem.input_memory_i.memory_wdata[62] ,
    \efabless_subsystem.input_memory_i.memory_wdata[61] ,
    \efabless_subsystem.input_memory_i.memory_wdata[60] ,
    \efabless_subsystem.input_memory_i.memory_wdata[59] ,
    \efabless_subsystem.input_memory_i.memory_wdata[58] ,
    \efabless_subsystem.input_memory_i.memory_wdata[57] ,
    \efabless_subsystem.input_memory_i.memory_wdata[56] ,
    \efabless_subsystem.input_memory_i.memory_wdata[55] ,
    \efabless_subsystem.input_memory_i.memory_wdata[54] ,
    \efabless_subsystem.input_memory_i.memory_wdata[53] ,
    \efabless_subsystem.input_memory_i.memory_wdata[52] ,
    \efabless_subsystem.input_memory_i.memory_wdata[51] ,
    \efabless_subsystem.input_memory_i.memory_wdata[50] ,
    \efabless_subsystem.input_memory_i.memory_wdata[49] ,
    \efabless_subsystem.input_memory_i.memory_wdata[48] ,
    \efabless_subsystem.input_memory_i.memory_wdata[47] ,
    \efabless_subsystem.input_memory_i.memory_wdata[46] ,
    \efabless_subsystem.input_memory_i.memory_wdata[45] ,
    \efabless_subsystem.input_memory_i.memory_wdata[44] ,
    \efabless_subsystem.input_memory_i.memory_wdata[43] ,
    \efabless_subsystem.input_memory_i.memory_wdata[42] ,
    \efabless_subsystem.input_memory_i.memory_wdata[41] ,
    \efabless_subsystem.input_memory_i.memory_wdata[40] ,
    \efabless_subsystem.input_memory_i.memory_wdata[39] ,
    \efabless_subsystem.input_memory_i.memory_wdata[38] ,
    \efabless_subsystem.input_memory_i.memory_wdata[37] ,
    \efabless_subsystem.input_memory_i.memory_wdata[36] ,
    \efabless_subsystem.input_memory_i.memory_wdata[35] ,
    \efabless_subsystem.input_memory_i.memory_wdata[34] ,
    \efabless_subsystem.input_memory_i.memory_wdata[33] ,
    \efabless_subsystem.input_memory_i.memory_wdata[32] ,
    \efabless_subsystem.input_memory_i.memory_wdata[31] ,
    \efabless_subsystem.input_memory_i.memory_wdata[30] ,
    \efabless_subsystem.input_memory_i.memory_wdata[29] ,
    \efabless_subsystem.input_memory_i.memory_wdata[28] ,
    \efabless_subsystem.input_memory_i.memory_wdata[27] ,
    \efabless_subsystem.input_memory_i.memory_wdata[26] ,
    \efabless_subsystem.input_memory_i.memory_wdata[25] ,
    \efabless_subsystem.input_memory_i.memory_wdata[24] ,
    \efabless_subsystem.input_memory_i.memory_wdata[23] ,
    \efabless_subsystem.input_memory_i.memory_wdata[22] ,
    \efabless_subsystem.input_memory_i.memory_wdata[21] ,
    \efabless_subsystem.input_memory_i.memory_wdata[20] ,
    \efabless_subsystem.input_memory_i.memory_wdata[19] ,
    \efabless_subsystem.input_memory_i.memory_wdata[18] ,
    \efabless_subsystem.input_memory_i.memory_wdata[17] ,
    \efabless_subsystem.input_memory_i.memory_wdata[16] ,
    \efabless_subsystem.input_memory_i.memory_wdata[15] ,
    \efabless_subsystem.input_memory_i.memory_wdata[14] ,
    \efabless_subsystem.input_memory_i.memory_wdata[13] ,
    \efabless_subsystem.input_memory_i.memory_wdata[12] ,
    \efabless_subsystem.input_memory_i.memory_wdata[11] ,
    \efabless_subsystem.input_memory_i.memory_wdata[10] ,
    \efabless_subsystem.input_memory_i.memory_wdata[9] ,
    \efabless_subsystem.input_memory_i.memory_wdata[8] ,
    \efabless_subsystem.input_memory_i.memory_wdata[7] ,
    \efabless_subsystem.input_memory_i.memory_wdata[6] ,
    \efabless_subsystem.input_memory_i.memory_wdata[5] ,
    \efabless_subsystem.input_memory_i.memory_wdata[4] ,
    \efabless_subsystem.input_memory_i.memory_wdata[3] ,
    \efabless_subsystem.input_memory_i.memory_wdata[2] ,
    \efabless_subsystem.input_memory_i.memory_wdata[1] ,
    \efabless_subsystem.input_memory_i.memory_wdata[0] }),
    .dout0({\efabless_subsystem.input_memory_i._009_ ,
    \efabless_subsystem.input_memory_i._008_ ,
    \efabless_subsystem.input_memory_i._007_ ,
    \efabless_subsystem.imem_rdata[196] ,
    \efabless_subsystem.imem_rdata[195] ,
    \efabless_subsystem.imem_rdata[194] ,
    \efabless_subsystem.imem_rdata[193] ,
    \efabless_subsystem.imem_rdata[192] ,
    \efabless_subsystem.imem_rdata[191] ,
    \efabless_subsystem.imem_rdata[190] ,
    \efabless_subsystem.imem_rdata[189] ,
    \efabless_subsystem.imem_rdata[188] ,
    \efabless_subsystem.imem_rdata[187] ,
    \efabless_subsystem.imem_rdata[186] ,
    \efabless_subsystem.imem_rdata[185] ,
    \efabless_subsystem.imem_rdata[184] ,
    \efabless_subsystem.imem_rdata[183] ,
    \efabless_subsystem.imem_rdata[182] ,
    \efabless_subsystem.imem_rdata[181] ,
    \efabless_subsystem.imem_rdata[180] ,
    \efabless_subsystem.imem_rdata[179] ,
    \efabless_subsystem.imem_rdata[178] ,
    \efabless_subsystem.imem_rdata[177] ,
    \efabless_subsystem.imem_rdata[176] ,
    \efabless_subsystem.imem_rdata[175] ,
    \efabless_subsystem.imem_rdata[174] ,
    \efabless_subsystem.imem_rdata[173] ,
    \efabless_subsystem.imem_rdata[172] ,
    \efabless_subsystem.imem_rdata[171] ,
    \efabless_subsystem.imem_rdata[170] ,
    \efabless_subsystem.imem_rdata[169] ,
    \efabless_subsystem.imem_rdata[168] ,
    \efabless_subsystem.imem_rdata[167] ,
    \efabless_subsystem.imem_rdata[166] ,
    \efabless_subsystem.imem_rdata[165] ,
    \efabless_subsystem.imem_rdata[164] ,
    \efabless_subsystem.imem_rdata[163] ,
    \efabless_subsystem.imem_rdata[162] ,
    \efabless_subsystem.imem_rdata[161] ,
    \efabless_subsystem.imem_rdata[160] ,
    \efabless_subsystem.imem_rdata[159] ,
    \efabless_subsystem.imem_rdata[158] ,
    \efabless_subsystem.imem_rdata[157] ,
    \efabless_subsystem.imem_rdata[156] ,
    \efabless_subsystem.imem_rdata[155] ,
    \efabless_subsystem.imem_rdata[154] ,
    \efabless_subsystem.imem_rdata[153] ,
    \efabless_subsystem.imem_rdata[152] ,
    \efabless_subsystem.imem_rdata[151] ,
    \efabless_subsystem.imem_rdata[150] ,
    \efabless_subsystem.imem_rdata[149] ,
    \efabless_subsystem.imem_rdata[148] ,
    \efabless_subsystem.imem_rdata[147] ,
    \efabless_subsystem.imem_rdata[146] ,
    \efabless_subsystem.imem_rdata[145] ,
    \efabless_subsystem.imem_rdata[144] ,
    \efabless_subsystem.imem_rdata[143] ,
    \efabless_subsystem.imem_rdata[142] ,
    \efabless_subsystem.imem_rdata[141] ,
    \efabless_subsystem.imem_rdata[140] ,
    \efabless_subsystem.imem_rdata[139] ,
    \efabless_subsystem.imem_rdata[138] ,
    \efabless_subsystem.imem_rdata[137] ,
    \efabless_subsystem.imem_rdata[136] ,
    \efabless_subsystem.imem_rdata[135] ,
    \efabless_subsystem.imem_rdata[134] ,
    \efabless_subsystem.imem_rdata[133] ,
    \efabless_subsystem.imem_rdata[132] ,
    \efabless_subsystem.imem_rdata[131] ,
    \efabless_subsystem.imem_rdata[130] ,
    \efabless_subsystem.imem_rdata[129] ,
    \efabless_subsystem.imem_rdata[128] ,
    \efabless_subsystem.imem_rdata[127] ,
    \efabless_subsystem.imem_rdata[126] ,
    \efabless_subsystem.imem_rdata[125] ,
    \efabless_subsystem.imem_rdata[124] ,
    \efabless_subsystem.imem_rdata[123] ,
    \efabless_subsystem.imem_rdata[122] ,
    \efabless_subsystem.imem_rdata[121] ,
    \efabless_subsystem.imem_rdata[120] ,
    \efabless_subsystem.imem_rdata[119] ,
    \efabless_subsystem.imem_rdata[118] ,
    \efabless_subsystem.imem_rdata[117] ,
    \efabless_subsystem.imem_rdata[116] ,
    \efabless_subsystem.imem_rdata[115] ,
    \efabless_subsystem.imem_rdata[114] ,
    \efabless_subsystem.imem_rdata[113] ,
    \efabless_subsystem.imem_rdata[112] ,
    \efabless_subsystem.imem_rdata[111] ,
    \efabless_subsystem.imem_rdata[110] ,
    \efabless_subsystem.imem_rdata[109] ,
    \efabless_subsystem.imem_rdata[108] ,
    \efabless_subsystem.imem_rdata[107] ,
    \efabless_subsystem.imem_rdata[106] ,
    \efabless_subsystem.imem_rdata[105] ,
    \efabless_subsystem.imem_rdata[104] ,
    \efabless_subsystem.imem_rdata[103] ,
    \efabless_subsystem.imem_rdata[102] ,
    \efabless_subsystem.imem_rdata[101] ,
    \efabless_subsystem.imem_rdata[100] ,
    \efabless_subsystem.imem_rdata[99] ,
    \efabless_subsystem.imem_rdata[98] ,
    \efabless_subsystem.imem_rdata[97] ,
    \efabless_subsystem.imem_rdata[96] ,
    \efabless_subsystem.imem_rdata[95] ,
    \efabless_subsystem.imem_rdata[94] ,
    \efabless_subsystem.imem_rdata[93] ,
    \efabless_subsystem.imem_rdata[92] ,
    \efabless_subsystem.imem_rdata[91] ,
    \efabless_subsystem.imem_rdata[90] ,
    \efabless_subsystem.imem_rdata[89] ,
    \efabless_subsystem.imem_rdata[88] ,
    \efabless_subsystem.imem_rdata[87] ,
    \efabless_subsystem.imem_rdata[86] ,
    \efabless_subsystem.imem_rdata[85] ,
    \efabless_subsystem.imem_rdata[84] ,
    \efabless_subsystem.imem_rdata[83] ,
    \efabless_subsystem.imem_rdata[82] ,
    \efabless_subsystem.imem_rdata[81] ,
    \efabless_subsystem.imem_rdata[80] ,
    \efabless_subsystem.imem_rdata[79] ,
    \efabless_subsystem.imem_rdata[78] ,
    \efabless_subsystem.imem_rdata[77] ,
    \efabless_subsystem.imem_rdata[76] ,
    \efabless_subsystem.imem_rdata[75] ,
    \efabless_subsystem.imem_rdata[74] ,
    \efabless_subsystem.imem_rdata[73] ,
    \efabless_subsystem.imem_rdata[72] ,
    \efabless_subsystem.imem_rdata[71] ,
    \efabless_subsystem.imem_rdata[70] ,
    \efabless_subsystem.imem_rdata[69] ,
    \efabless_subsystem.imem_rdata[68] ,
    \efabless_subsystem.imem_rdata[67] ,
    \efabless_subsystem.imem_rdata[66] ,
    \efabless_subsystem.imem_rdata[65] ,
    \efabless_subsystem.imem_rdata[64] ,
    \efabless_subsystem.imem_rdata[63] ,
    \efabless_subsystem.imem_rdata[62] ,
    \efabless_subsystem.imem_rdata[61] ,
    \efabless_subsystem.imem_rdata[60] ,
    \efabless_subsystem.imem_rdata[59] ,
    \efabless_subsystem.imem_rdata[58] ,
    \efabless_subsystem.imem_rdata[57] ,
    \efabless_subsystem.imem_rdata[56] ,
    \efabless_subsystem.imem_rdata[55] ,
    \efabless_subsystem.imem_rdata[54] ,
    \efabless_subsystem.imem_rdata[53] ,
    \efabless_subsystem.imem_rdata[52] ,
    \efabless_subsystem.imem_rdata[51] ,
    \efabless_subsystem.imem_rdata[50] ,
    \efabless_subsystem.imem_rdata[49] ,
    \efabless_subsystem.imem_rdata[48] ,
    \efabless_subsystem.imem_rdata[47] ,
    \efabless_subsystem.imem_rdata[46] ,
    \efabless_subsystem.imem_rdata[45] ,
    \efabless_subsystem.imem_rdata[44] ,
    \efabless_subsystem.imem_rdata[43] ,
    \efabless_subsystem.imem_rdata[42] ,
    \efabless_subsystem.imem_rdata[41] ,
    \efabless_subsystem.imem_rdata[40] ,
    \efabless_subsystem.imem_rdata[39] ,
    \efabless_subsystem.imem_rdata[38] ,
    \efabless_subsystem.imem_rdata[37] ,
    \efabless_subsystem.imem_rdata[36] ,
    \efabless_subsystem.imem_rdata[35] ,
    \efabless_subsystem.imem_rdata[34] ,
    \efabless_subsystem.imem_rdata[33] ,
    \efabless_subsystem.imem_rdata[32] ,
    \efabless_subsystem.imem_rdata[31] ,
    \efabless_subsystem.imem_rdata[30] ,
    \efabless_subsystem.imem_rdata[29] ,
    \efabless_subsystem.imem_rdata[28] ,
    \efabless_subsystem.imem_rdata[27] ,
    \efabless_subsystem.imem_rdata[26] ,
    \efabless_subsystem.imem_rdata[25] ,
    \efabless_subsystem.imem_rdata[24] ,
    \efabless_subsystem.imem_rdata[23] ,
    \efabless_subsystem.imem_rdata[22] ,
    \efabless_subsystem.imem_rdata[21] ,
    \efabless_subsystem.imem_rdata[20] ,
    \efabless_subsystem.imem_rdata[19] ,
    \efabless_subsystem.imem_rdata[18] ,
    \efabless_subsystem.imem_rdata[17] ,
    \efabless_subsystem.imem_rdata[16] ,
    \efabless_subsystem.imem_rdata[15] ,
    \efabless_subsystem.imem_rdata[14] ,
    \efabless_subsystem.imem_rdata[13] ,
    \efabless_subsystem.imem_rdata[12] ,
    \efabless_subsystem.imem_rdata[11] ,
    \efabless_subsystem.imem_rdata[10] ,
    \efabless_subsystem.imem_rdata[9] ,
    \efabless_subsystem.imem_rdata[8] ,
    \efabless_subsystem.imem_rdata[7] ,
    \efabless_subsystem.imem_rdata[6] ,
    \efabless_subsystem.imem_rdata[5] ,
    \efabless_subsystem.imem_rdata[4] ,
    \efabless_subsystem.imem_rdata[3] ,
    \efabless_subsystem.imem_rdata[2] ,
    \efabless_subsystem.imem_rdata[1] ,
    \efabless_subsystem.imem_rdata[0] }),
    .dout1({\efabless_subsystem.input_memory_i._006_ ,
    \efabless_subsystem.input_memory_i._005_ ,
    \efabless_subsystem.input_memory_i._004_ ,
    \efabless_subsystem.core_stat_data_valid ,
    \efabless_subsystem.compute_core_i.i_array_shftsgn[3] ,
    \efabless_subsystem.compute_core_i.i_array_shftsgn[2] ,
    \efabless_subsystem.compute_core_i.i_array_shftsgn[1] ,
    \efabless_subsystem.compute_core_i.i_array_shftsgn[0] ,
    \efabless_subsystem.compute_core_i.i_weight[127] ,
    \efabless_subsystem.compute_core_i.i_weight[126] ,
    \efabless_subsystem.compute_core_i.i_weight[125] ,
    \efabless_subsystem.compute_core_i.i_weight[124] ,
    \efabless_subsystem.compute_core_i.i_weight[123] ,
    \efabless_subsystem.compute_core_i.i_weight[122] ,
    \efabless_subsystem.compute_core_i.i_weight[121] ,
    \efabless_subsystem.compute_core_i.i_weight[120] ,
    \efabless_subsystem.compute_core_i.i_weight[119] ,
    \efabless_subsystem.compute_core_i.i_weight[118] ,
    \efabless_subsystem.compute_core_i.i_weight[117] ,
    \efabless_subsystem.compute_core_i.i_weight[116] ,
    \efabless_subsystem.compute_core_i.i_weight[115] ,
    \efabless_subsystem.compute_core_i.i_weight[114] ,
    \efabless_subsystem.compute_core_i.i_weight[113] ,
    \efabless_subsystem.compute_core_i.i_weight[112] ,
    \efabless_subsystem.compute_core_i.i_weight[111] ,
    \efabless_subsystem.compute_core_i.i_weight[110] ,
    \efabless_subsystem.compute_core_i.i_weight[109] ,
    \efabless_subsystem.compute_core_i.i_weight[108] ,
    \efabless_subsystem.compute_core_i.i_weight[107] ,
    \efabless_subsystem.compute_core_i.i_weight[106] ,
    \efabless_subsystem.compute_core_i.i_weight[105] ,
    \efabless_subsystem.compute_core_i.i_weight[104] ,
    \efabless_subsystem.compute_core_i.i_weight[103] ,
    \efabless_subsystem.compute_core_i.i_weight[102] ,
    \efabless_subsystem.compute_core_i.i_weight[101] ,
    \efabless_subsystem.compute_core_i.i_weight[100] ,
    \efabless_subsystem.compute_core_i.i_weight[99] ,
    \efabless_subsystem.compute_core_i.i_weight[98] ,
    \efabless_subsystem.compute_core_i.i_weight[97] ,
    \efabless_subsystem.compute_core_i.i_weight[96] ,
    \efabless_subsystem.compute_core_i.i_weight[95] ,
    \efabless_subsystem.compute_core_i.i_weight[94] ,
    \efabless_subsystem.compute_core_i.i_weight[93] ,
    \efabless_subsystem.compute_core_i.i_weight[92] ,
    \efabless_subsystem.compute_core_i.i_weight[91] ,
    \efabless_subsystem.compute_core_i.i_weight[90] ,
    \efabless_subsystem.compute_core_i.i_weight[89] ,
    \efabless_subsystem.compute_core_i.i_weight[88] ,
    \efabless_subsystem.compute_core_i.i_weight[87] ,
    \efabless_subsystem.compute_core_i.i_weight[86] ,
    \efabless_subsystem.compute_core_i.i_weight[85] ,
    \efabless_subsystem.compute_core_i.i_weight[84] ,
    \efabless_subsystem.compute_core_i.i_weight[83] ,
    \efabless_subsystem.compute_core_i.i_weight[82] ,
    \efabless_subsystem.compute_core_i.i_weight[81] ,
    \efabless_subsystem.compute_core_i.i_weight[80] ,
    \efabless_subsystem.compute_core_i.i_weight[79] ,
    \efabless_subsystem.compute_core_i.i_weight[78] ,
    \efabless_subsystem.compute_core_i.i_weight[77] ,
    \efabless_subsystem.compute_core_i.i_weight[76] ,
    \efabless_subsystem.compute_core_i.i_weight[75] ,
    \efabless_subsystem.compute_core_i.i_weight[74] ,
    \efabless_subsystem.compute_core_i.i_weight[73] ,
    \efabless_subsystem.compute_core_i.i_weight[72] ,
    \efabless_subsystem.compute_core_i.i_weight[71] ,
    \efabless_subsystem.compute_core_i.i_weight[70] ,
    \efabless_subsystem.compute_core_i.i_weight[69] ,
    \efabless_subsystem.compute_core_i.i_weight[68] ,
    \efabless_subsystem.compute_core_i.i_weight[67] ,
    \efabless_subsystem.compute_core_i.i_weight[66] ,
    \efabless_subsystem.compute_core_i.i_weight[65] ,
    \efabless_subsystem.compute_core_i.i_weight[64] ,
    \efabless_subsystem.compute_core_i.i_weight[63] ,
    \efabless_subsystem.compute_core_i.i_weight[62] ,
    \efabless_subsystem.compute_core_i.i_weight[61] ,
    \efabless_subsystem.compute_core_i.i_weight[60] ,
    \efabless_subsystem.compute_core_i.i_weight[59] ,
    \efabless_subsystem.compute_core_i.i_weight[58] ,
    \efabless_subsystem.compute_core_i.i_weight[57] ,
    \efabless_subsystem.compute_core_i.i_weight[56] ,
    \efabless_subsystem.compute_core_i.i_weight[55] ,
    \efabless_subsystem.compute_core_i.i_weight[54] ,
    \efabless_subsystem.compute_core_i.i_weight[53] ,
    \efabless_subsystem.compute_core_i.i_weight[52] ,
    \efabless_subsystem.compute_core_i.i_weight[51] ,
    \efabless_subsystem.compute_core_i.i_weight[50] ,
    \efabless_subsystem.compute_core_i.i_weight[49] ,
    \efabless_subsystem.compute_core_i.i_weight[48] ,
    \efabless_subsystem.compute_core_i.i_weight[47] ,
    \efabless_subsystem.compute_core_i.i_weight[46] ,
    \efabless_subsystem.compute_core_i.i_weight[45] ,
    \efabless_subsystem.compute_core_i.i_weight[44] ,
    \efabless_subsystem.compute_core_i.i_weight[43] ,
    \efabless_subsystem.compute_core_i.i_weight[42] ,
    \efabless_subsystem.compute_core_i.i_weight[41] ,
    \efabless_subsystem.compute_core_i.i_weight[40] ,
    \efabless_subsystem.compute_core_i.i_weight[39] ,
    \efabless_subsystem.compute_core_i.i_weight[38] ,
    \efabless_subsystem.compute_core_i.i_weight[37] ,
    \efabless_subsystem.compute_core_i.i_weight[36] ,
    \efabless_subsystem.compute_core_i.i_weight[35] ,
    \efabless_subsystem.compute_core_i.i_weight[34] ,
    \efabless_subsystem.compute_core_i.i_weight[33] ,
    \efabless_subsystem.compute_core_i.i_weight[32] ,
    \efabless_subsystem.compute_core_i.i_weight[31] ,
    \efabless_subsystem.compute_core_i.i_weight[30] ,
    \efabless_subsystem.compute_core_i.i_weight[29] ,
    \efabless_subsystem.compute_core_i.i_weight[28] ,
    \efabless_subsystem.compute_core_i.i_weight[27] ,
    \efabless_subsystem.compute_core_i.i_weight[26] ,
    \efabless_subsystem.compute_core_i.i_weight[25] ,
    \efabless_subsystem.compute_core_i.i_weight[24] ,
    \efabless_subsystem.compute_core_i.i_weight[23] ,
    \efabless_subsystem.compute_core_i.i_weight[22] ,
    \efabless_subsystem.compute_core_i.i_weight[21] ,
    \efabless_subsystem.compute_core_i.i_weight[20] ,
    \efabless_subsystem.compute_core_i.i_weight[19] ,
    \efabless_subsystem.compute_core_i.i_weight[18] ,
    \efabless_subsystem.compute_core_i.i_weight[17] ,
    \efabless_subsystem.compute_core_i.i_weight[16] ,
    \efabless_subsystem.compute_core_i.i_weight[15] ,
    \efabless_subsystem.compute_core_i.i_weight[14] ,
    \efabless_subsystem.compute_core_i.i_weight[13] ,
    \efabless_subsystem.compute_core_i.i_weight[12] ,
    \efabless_subsystem.compute_core_i.i_weight[11] ,
    \efabless_subsystem.compute_core_i.i_weight[10] ,
    \efabless_subsystem.compute_core_i.i_weight[9] ,
    \efabless_subsystem.compute_core_i.i_weight[8] ,
    \efabless_subsystem.compute_core_i.i_weight[7] ,
    \efabless_subsystem.compute_core_i.i_weight[6] ,
    \efabless_subsystem.compute_core_i.i_weight[5] ,
    \efabless_subsystem.compute_core_i.i_weight[4] ,
    \efabless_subsystem.compute_core_i.i_weight[3] ,
    \efabless_subsystem.compute_core_i.i_weight[2] ,
    \efabless_subsystem.compute_core_i.i_weight[1] ,
    \efabless_subsystem.compute_core_i.i_weight[0] ,
    \efabless_subsystem.compute_core_i.i_fmap[63] ,
    \efabless_subsystem.compute_core_i.i_fmap[62] ,
    \efabless_subsystem.compute_core_i.i_fmap[61] ,
    \efabless_subsystem.compute_core_i.i_fmap[60] ,
    \efabless_subsystem.compute_core_i.i_fmap[59] ,
    \efabless_subsystem.compute_core_i.i_fmap[58] ,
    \efabless_subsystem.compute_core_i.i_fmap[57] ,
    \efabless_subsystem.compute_core_i.i_fmap[56] ,
    \efabless_subsystem.compute_core_i.i_fmap[55] ,
    \efabless_subsystem.compute_core_i.i_fmap[54] ,
    \efabless_subsystem.compute_core_i.i_fmap[53] ,
    \efabless_subsystem.compute_core_i.i_fmap[52] ,
    \efabless_subsystem.compute_core_i.i_fmap[51] ,
    \efabless_subsystem.compute_core_i.i_fmap[50] ,
    \efabless_subsystem.compute_core_i.i_fmap[49] ,
    \efabless_subsystem.compute_core_i.i_fmap[48] ,
    \efabless_subsystem.compute_core_i.i_fmap[47] ,
    \efabless_subsystem.compute_core_i.i_fmap[46] ,
    \efabless_subsystem.compute_core_i.i_fmap[45] ,
    \efabless_subsystem.compute_core_i.i_fmap[44] ,
    \efabless_subsystem.compute_core_i.i_fmap[43] ,
    \efabless_subsystem.compute_core_i.i_fmap[42] ,
    \efabless_subsystem.compute_core_i.i_fmap[41] ,
    \efabless_subsystem.compute_core_i.i_fmap[40] ,
    \efabless_subsystem.compute_core_i.i_fmap[39] ,
    \efabless_subsystem.compute_core_i.i_fmap[38] ,
    \efabless_subsystem.compute_core_i.i_fmap[37] ,
    \efabless_subsystem.compute_core_i.i_fmap[36] ,
    \efabless_subsystem.compute_core_i.i_fmap[35] ,
    \efabless_subsystem.compute_core_i.i_fmap[34] ,
    \efabless_subsystem.compute_core_i.i_fmap[33] ,
    \efabless_subsystem.compute_core_i.i_fmap[32] ,
    \efabless_subsystem.compute_core_i.i_fmap[31] ,
    \efabless_subsystem.compute_core_i.i_fmap[30] ,
    \efabless_subsystem.compute_core_i.i_fmap[29] ,
    \efabless_subsystem.compute_core_i.i_fmap[28] ,
    \efabless_subsystem.compute_core_i.i_fmap[27] ,
    \efabless_subsystem.compute_core_i.i_fmap[26] ,
    \efabless_subsystem.compute_core_i.i_fmap[25] ,
    \efabless_subsystem.compute_core_i.i_fmap[24] ,
    \efabless_subsystem.compute_core_i.i_fmap[23] ,
    \efabless_subsystem.compute_core_i.i_fmap[22] ,
    \efabless_subsystem.compute_core_i.i_fmap[21] ,
    \efabless_subsystem.compute_core_i.i_fmap[20] ,
    \efabless_subsystem.compute_core_i.i_fmap[19] ,
    \efabless_subsystem.compute_core_i.i_fmap[18] ,
    \efabless_subsystem.compute_core_i.i_fmap[17] ,
    \efabless_subsystem.compute_core_i.i_fmap[16] ,
    \efabless_subsystem.compute_core_i.i_fmap[15] ,
    \efabless_subsystem.compute_core_i.i_fmap[14] ,
    \efabless_subsystem.compute_core_i.i_fmap[13] ,
    \efabless_subsystem.compute_core_i.i_fmap[12] ,
    \efabless_subsystem.compute_core_i.i_fmap[11] ,
    \efabless_subsystem.compute_core_i.i_fmap[10] ,
    \efabless_subsystem.compute_core_i.i_fmap[9] ,
    \efabless_subsystem.compute_core_i.i_fmap[8] ,
    \efabless_subsystem.compute_core_i.i_fmap[7] ,
    \efabless_subsystem.compute_core_i.i_fmap[6] ,
    \efabless_subsystem.compute_core_i.i_fmap[5] ,
    \efabless_subsystem.compute_core_i.i_fmap[4] ,
    \efabless_subsystem.compute_core_i.i_fmap[3] ,
    \efabless_subsystem.compute_core_i.i_fmap[2] ,
    \efabless_subsystem.compute_core_i.i_fmap[1] ,
    \efabless_subsystem.compute_core_i.i_fmap[0] }),
    .wmask0({\efabless_subsystem.input_memory_i.memory_wmask[24] ,
    \efabless_subsystem.input_memory_i.memory_wmask[23] ,
    \efabless_subsystem.input_memory_i.memory_wmask[22] ,
    \efabless_subsystem.input_memory_i.memory_wmask[21] ,
    \efabless_subsystem.input_memory_i.memory_wmask[20] ,
    \efabless_subsystem.input_memory_i.memory_wmask[19] ,
    \efabless_subsystem.input_memory_i.memory_wmask[18] ,
    \efabless_subsystem.input_memory_i.memory_wmask[17] ,
    \efabless_subsystem.input_memory_i.memory_wmask[16] ,
    \efabless_subsystem.input_memory_i.memory_wmask[15] ,
    \efabless_subsystem.input_memory_i.memory_wmask[14] ,
    \efabless_subsystem.input_memory_i.memory_wmask[13] ,
    \efabless_subsystem.input_memory_i.memory_wmask[12] ,
    \efabless_subsystem.input_memory_i.memory_wmask[11] ,
    \efabless_subsystem.input_memory_i.memory_wmask[10] ,
    \efabless_subsystem.input_memory_i.memory_wmask[9] ,
    \efabless_subsystem.input_memory_i.memory_wmask[8] ,
    \efabless_subsystem.input_memory_i.memory_wmask[7] ,
    \efabless_subsystem.input_memory_i.memory_wmask[6] ,
    \efabless_subsystem.input_memory_i.memory_wmask[5] ,
    \efabless_subsystem.input_memory_i.memory_wmask[4] ,
    \efabless_subsystem.input_memory_i.memory_wmask[3] ,
    \efabless_subsystem.input_memory_i.memory_wmask[2] ,
    \efabless_subsystem.input_memory_i.memory_wmask[1] ,
    \efabless_subsystem.input_memory_i.memory_wmask[0] }));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g1._1_  (.A0(\efabless_subsystem.imem_wdata[196] ),
    .A1(\efabless_subsystem._199_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[196] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g10._1_  (.A0(\efabless_subsystem.imem_wdata[187] ),
    .A1(\efabless_subsystem._190_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[187] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g100._1_  (.A0(\efabless_subsystem.imem_wdata[97] ),
    .A1(\efabless_subsystem._100_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g100._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g100._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g100._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[97] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g101._1_  (.A0(\efabless_subsystem.imem_wdata[96] ),
    .A1(\efabless_subsystem._099_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g101._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g101._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g101._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[96] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g102._1_  (.A0(\efabless_subsystem.imem_wdata[95] ),
    .A1(\efabless_subsystem._098_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g102._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g102._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g102._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[95] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g103._1_  (.A0(\efabless_subsystem.imem_wdata[94] ),
    .A1(\efabless_subsystem._097_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g103._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g103._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g103._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[94] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g104._1_  (.A0(\efabless_subsystem.imem_wdata[93] ),
    .A1(\efabless_subsystem._096_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g104._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g104._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g104._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[93] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g105._1_  (.A0(\efabless_subsystem.imem_wdata[92] ),
    .A1(\efabless_subsystem._095_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g105._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g105._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g105._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[92] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g106._1_  (.A0(\efabless_subsystem.imem_wdata[91] ),
    .A1(\efabless_subsystem._094_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g106._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g106._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g106._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[91] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g107._1_  (.A0(\efabless_subsystem.imem_wdata[90] ),
    .A1(\efabless_subsystem._093_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g107._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g107._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g107._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[90] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g108._1_  (.A0(\efabless_subsystem.imem_wdata[89] ),
    .A1(\efabless_subsystem._092_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g108._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g108._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g108._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[89] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g109._1_  (.A0(\efabless_subsystem.imem_wdata[88] ),
    .A1(\efabless_subsystem._091_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g109._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g109._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g109._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[88] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g11._1_  (.A0(\efabless_subsystem.imem_wdata[186] ),
    .A1(\efabless_subsystem._189_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[186] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g110._1_  (.A0(\efabless_subsystem.imem_wdata[87] ),
    .A1(\efabless_subsystem._090_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g110._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g110._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g110._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[87] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g111._1_  (.A0(\efabless_subsystem.imem_wdata[86] ),
    .A1(\efabless_subsystem._089_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g111._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g111._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g111._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[86] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g112._1_  (.A0(\efabless_subsystem.imem_wdata[85] ),
    .A1(\efabless_subsystem._088_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g112._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g112._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g112._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[85] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g113._1_  (.A0(\efabless_subsystem.imem_wdata[84] ),
    .A1(\efabless_subsystem._087_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g113._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g113._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g113._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[84] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g114._1_  (.A0(\efabless_subsystem.imem_wdata[83] ),
    .A1(\efabless_subsystem._086_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g114._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g114._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g114._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[83] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g115._1_  (.A0(\efabless_subsystem.imem_wdata[82] ),
    .A1(\efabless_subsystem._085_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g115._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g115._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g115._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[82] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g116._1_  (.A0(\efabless_subsystem.imem_wdata[81] ),
    .A1(\efabless_subsystem._084_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g116._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g116._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g116._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[81] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g117._1_  (.A0(\efabless_subsystem.imem_wdata[80] ),
    .A1(\efabless_subsystem._083_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g117._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g117._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g117._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[80] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g118._1_  (.A0(\efabless_subsystem.imem_wdata[79] ),
    .A1(\efabless_subsystem._082_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g118._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g118._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g118._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[79] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g119._1_  (.A0(\efabless_subsystem.imem_wdata[78] ),
    .A1(\efabless_subsystem._081_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g119._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g119._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g119._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[78] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g12._1_  (.A0(\efabless_subsystem.imem_wdata[185] ),
    .A1(\efabless_subsystem._188_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[185] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g120._1_  (.A0(\efabless_subsystem.imem_wdata[77] ),
    .A1(\efabless_subsystem._080_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g120._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g120._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g120._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[77] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g121._1_  (.A0(\efabless_subsystem.imem_wdata[76] ),
    .A1(\efabless_subsystem._079_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g121._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g121._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g121._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[76] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g122._1_  (.A0(\efabless_subsystem.imem_wdata[75] ),
    .A1(\efabless_subsystem._078_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g122._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g122._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g122._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[75] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g123._1_  (.A0(\efabless_subsystem.imem_wdata[74] ),
    .A1(\efabless_subsystem._077_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g123._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g123._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g123._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[74] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g124._1_  (.A0(\efabless_subsystem.imem_wdata[73] ),
    .A1(\efabless_subsystem._076_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g124._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g124._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g124._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[73] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g125._1_  (.A0(\efabless_subsystem.imem_wdata[72] ),
    .A1(\efabless_subsystem._075_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g125._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g125._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g125._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[72] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g126._1_  (.A0(\efabless_subsystem.imem_wdata[71] ),
    .A1(\efabless_subsystem._074_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g126._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g126._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g126._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[71] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g127._1_  (.A0(\efabless_subsystem.imem_wdata[70] ),
    .A1(\efabless_subsystem._073_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g127._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g127._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g127._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[70] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g128._1_  (.A0(\efabless_subsystem.imem_wdata[69] ),
    .A1(\efabless_subsystem._072_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g128._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g128._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g128._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[69] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g129._1_  (.A0(\efabless_subsystem.imem_wdata[68] ),
    .A1(\efabless_subsystem._071_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g129._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g129._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g129._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[68] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g13._1_  (.A0(\efabless_subsystem.imem_wdata[184] ),
    .A1(\efabless_subsystem._187_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g13._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[184] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g130._1_  (.A0(\efabless_subsystem.imem_wdata[67] ),
    .A1(\efabless_subsystem._070_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g130._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g130._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g130._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[67] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g131._1_  (.A0(\efabless_subsystem.imem_wdata[66] ),
    .A1(\efabless_subsystem._069_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g131._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g131._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g131._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[66] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g132._1_  (.A0(\efabless_subsystem.imem_wdata[65] ),
    .A1(\efabless_subsystem._068_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g132._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g132._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g132._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[65] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g133._1_  (.A0(\efabless_subsystem.imem_wdata[64] ),
    .A1(\efabless_subsystem._067_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g133._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g133._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g133._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[64] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g134._1_  (.A0(\efabless_subsystem.imem_wdata[63] ),
    .A1(\efabless_subsystem._066_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g134._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g134._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g134._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[63] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g135._1_  (.A0(\efabless_subsystem.imem_wdata[62] ),
    .A1(\efabless_subsystem._065_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g135._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g135._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g135._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[62] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g136._1_  (.A0(\efabless_subsystem.imem_wdata[61] ),
    .A1(\efabless_subsystem._064_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g136._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g136._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g136._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[61] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g137._1_  (.A0(\efabless_subsystem.imem_wdata[60] ),
    .A1(\efabless_subsystem._063_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g137._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g137._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g137._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[60] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g138._1_  (.A0(\efabless_subsystem.imem_wdata[59] ),
    .A1(\efabless_subsystem._062_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g138._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g138._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g138._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[59] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g139._1_  (.A0(\efabless_subsystem.imem_wdata[58] ),
    .A1(\efabless_subsystem._061_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g139._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g139._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g139._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[58] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g14._1_  (.A0(\efabless_subsystem.imem_wdata[183] ),
    .A1(\efabless_subsystem._186_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g14._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[183] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g140._1_  (.A0(\efabless_subsystem.imem_wdata[57] ),
    .A1(\efabless_subsystem._060_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g140._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g140._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g140._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[57] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g141._1_  (.A0(\efabless_subsystem.imem_wdata[56] ),
    .A1(\efabless_subsystem._059_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g141._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g141._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g141._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[56] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g142._1_  (.A0(\efabless_subsystem.imem_wdata[55] ),
    .A1(\efabless_subsystem._058_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g142._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g142._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g142._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[55] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g143._1_  (.A0(\efabless_subsystem.imem_wdata[54] ),
    .A1(\efabless_subsystem._057_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g143._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g143._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g143._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[54] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g144._1_  (.A0(\efabless_subsystem.imem_wdata[53] ),
    .A1(\efabless_subsystem._056_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g144._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g144._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g144._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[53] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g145._1_  (.A0(\efabless_subsystem.imem_wdata[52] ),
    .A1(\efabless_subsystem._055_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g145._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g145._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g145._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[52] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g146._1_  (.A0(\efabless_subsystem.imem_wdata[51] ),
    .A1(\efabless_subsystem._054_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g146._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g146._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g146._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[51] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g147._1_  (.A0(\efabless_subsystem.imem_wdata[50] ),
    .A1(\efabless_subsystem._053_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g147._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g147._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g147._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[50] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g148._1_  (.A0(\efabless_subsystem.imem_wdata[49] ),
    .A1(\efabless_subsystem._052_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g148._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g148._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g148._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[49] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g149._1_  (.A0(\efabless_subsystem.imem_wdata[48] ),
    .A1(\efabless_subsystem._051_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g149._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g149._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g149._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[48] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g15._1_  (.A0(\efabless_subsystem.imem_wdata[182] ),
    .A1(\efabless_subsystem._185_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g15._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[182] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g150._1_  (.A0(\efabless_subsystem.imem_wdata[47] ),
    .A1(\efabless_subsystem._050_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g150._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g150._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g150._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[47] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g151._1_  (.A0(\efabless_subsystem.imem_wdata[46] ),
    .A1(\efabless_subsystem._049_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g151._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g151._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g151._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[46] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g152._1_  (.A0(\efabless_subsystem.imem_wdata[45] ),
    .A1(\efabless_subsystem._048_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g152._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g152._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g152._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[45] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g153._1_  (.A0(\efabless_subsystem.imem_wdata[44] ),
    .A1(\efabless_subsystem._047_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g153._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g153._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g153._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[44] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g154._1_  (.A0(\efabless_subsystem.imem_wdata[43] ),
    .A1(\efabless_subsystem._046_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g154._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g154._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g154._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[43] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g155._1_  (.A0(\efabless_subsystem.imem_wdata[42] ),
    .A1(\efabless_subsystem._045_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g155._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g155._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g155._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[42] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g156._1_  (.A0(\efabless_subsystem.imem_wdata[41] ),
    .A1(\efabless_subsystem._044_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g156._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g156._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g156._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[41] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g157._1_  (.A0(\efabless_subsystem.imem_wdata[40] ),
    .A1(\efabless_subsystem._043_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g157._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g157._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g157._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[40] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g158._1_  (.A0(\efabless_subsystem.imem_wdata[39] ),
    .A1(\efabless_subsystem._042_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g158._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g158._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g158._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[39] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g159._1_  (.A0(\efabless_subsystem.imem_wdata[38] ),
    .A1(\efabless_subsystem._041_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g159._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g159._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g159._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[38] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g16._1_  (.A0(\efabless_subsystem.imem_wdata[181] ),
    .A1(\efabless_subsystem._184_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g16._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[181] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g160._1_  (.A0(\efabless_subsystem.imem_wdata[37] ),
    .A1(\efabless_subsystem._040_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g160._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g160._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g160._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[37] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g161._1_  (.A0(\efabless_subsystem.imem_wdata[36] ),
    .A1(\efabless_subsystem._039_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g161._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g161._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g161._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[36] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g162._1_  (.A0(\efabless_subsystem.imem_wdata[35] ),
    .A1(\efabless_subsystem._038_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g162._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g162._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g162._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[35] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g163._1_  (.A0(\efabless_subsystem.imem_wdata[34] ),
    .A1(\efabless_subsystem._037_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g163._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g163._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g163._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[34] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g164._1_  (.A0(\efabless_subsystem.imem_wdata[33] ),
    .A1(\efabless_subsystem._036_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g164._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g164._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g164._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[33] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g165._1_  (.A0(\efabless_subsystem.imem_wdata[32] ),
    .A1(\efabless_subsystem._035_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g165._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g165._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g165._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[32] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g166._1_  (.A0(\efabless_subsystem.imem_wdata[31] ),
    .A1(\efabless_subsystem._034_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g166._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g166._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g166._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[31] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g167._1_  (.A0(\efabless_subsystem.imem_wdata[30] ),
    .A1(\efabless_subsystem._033_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g167._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g167._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g167._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[30] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g168._1_  (.A0(\efabless_subsystem.imem_wdata[29] ),
    .A1(\efabless_subsystem._032_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g168._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g168._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g168._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[29] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g169._1_  (.A0(\efabless_subsystem.imem_wdata[28] ),
    .A1(\efabless_subsystem._031_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g169._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g169._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g169._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[28] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g17._1_  (.A0(\efabless_subsystem.imem_wdata[180] ),
    .A1(\efabless_subsystem._183_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g17._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g17._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g17._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[180] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g170._1_  (.A0(\efabless_subsystem.imem_wdata[27] ),
    .A1(\efabless_subsystem._030_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g170._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g170._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g170._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[27] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g171._1_  (.A0(\efabless_subsystem.imem_wdata[26] ),
    .A1(\efabless_subsystem._029_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g171._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g171._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g171._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[26] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g172._1_  (.A0(\efabless_subsystem.imem_wdata[25] ),
    .A1(\efabless_subsystem._028_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g172._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g172._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g172._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[25] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g173._1_  (.A0(\efabless_subsystem.imem_wdata[24] ),
    .A1(\efabless_subsystem._027_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g173._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g173._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g173._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[24] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g174._1_  (.A0(\efabless_subsystem.imem_wdata[23] ),
    .A1(\efabless_subsystem._026_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g174._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g174._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g174._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[23] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g175._1_  (.A0(\efabless_subsystem.imem_wdata[22] ),
    .A1(\efabless_subsystem._025_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g175._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g175._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g175._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[22] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g176._1_  (.A0(\efabless_subsystem.imem_wdata[21] ),
    .A1(\efabless_subsystem._024_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g176._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g176._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g176._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[21] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g177._1_  (.A0(\efabless_subsystem.imem_wdata[20] ),
    .A1(\efabless_subsystem._023_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g177._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g177._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g177._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[20] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g178._1_  (.A0(\efabless_subsystem.imem_wdata[19] ),
    .A1(\efabless_subsystem._022_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g178._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g178._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g178._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[19] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g179._1_  (.A0(\efabless_subsystem.imem_wdata[18] ),
    .A1(\efabless_subsystem._021_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g179._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g179._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g179._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[18] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g18._1_  (.A0(\efabless_subsystem.imem_wdata[179] ),
    .A1(\efabless_subsystem._182_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g18._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g18._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g18._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[179] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g180._1_  (.A0(\efabless_subsystem.imem_wdata[17] ),
    .A1(\efabless_subsystem._020_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g180._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g180._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g180._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[17] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g181._1_  (.A0(\efabless_subsystem.imem_wdata[16] ),
    .A1(\efabless_subsystem._019_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g181._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g181._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g181._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[16] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g182._1_  (.A0(\efabless_subsystem.imem_wdata[15] ),
    .A1(\efabless_subsystem._018_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g182._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g182._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g182._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[15] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g183._1_  (.A0(\efabless_subsystem.imem_wdata[14] ),
    .A1(\efabless_subsystem._017_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g183._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g183._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g183._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[14] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g184._1_  (.A0(\efabless_subsystem.imem_wdata[13] ),
    .A1(\efabless_subsystem._016_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g184._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g184._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g184._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[13] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g185._1_  (.A0(\efabless_subsystem.imem_wdata[12] ),
    .A1(\efabless_subsystem._015_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g185._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g185._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g185._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[12] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g186._1_  (.A0(\efabless_subsystem.imem_wdata[11] ),
    .A1(\efabless_subsystem._014_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g186._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g186._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g186._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[11] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g187._1_  (.A0(\efabless_subsystem.imem_wdata[10] ),
    .A1(\efabless_subsystem._013_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g187._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g187._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g187._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[10] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g188._1_  (.A0(\efabless_subsystem.imem_wdata[9] ),
    .A1(\efabless_subsystem._012_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g188._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g188._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g188._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[9] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g189._1_  (.A0(\efabless_subsystem.imem_wdata[8] ),
    .A1(\efabless_subsystem._011_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g189._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g189._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g189._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[8] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g19._1_  (.A0(\efabless_subsystem.imem_wdata[178] ),
    .A1(\efabless_subsystem._181_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g19._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g19._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g19._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[178] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g190._1_  (.A0(\efabless_subsystem.imem_wdata[7] ),
    .A1(\efabless_subsystem._010_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g190._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g190._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g190._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[7] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g191._1_  (.A0(\efabless_subsystem.imem_wdata[6] ),
    .A1(\efabless_subsystem._009_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g191._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g191._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g191._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[6] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g192._1_  (.A0(\efabless_subsystem.imem_wdata[5] ),
    .A1(\efabless_subsystem._008_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g192._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g192._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g192._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[5] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g193._1_  (.A0(\efabless_subsystem.imem_wdata[4] ),
    .A1(\efabless_subsystem._007_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g193._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g193._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g193._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g194._1_  (.A0(\efabless_subsystem.imem_wdata[3] ),
    .A1(\efabless_subsystem._006_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g194._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g194._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g194._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g195._1_  (.A0(\efabless_subsystem.imem_wdata[2] ),
    .A1(\efabless_subsystem._005_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g195._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g195._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g195._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g196._1_  (.A0(\efabless_subsystem.imem_wdata[1] ),
    .A1(\efabless_subsystem._004_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g196._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g196._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g196._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g197._1_  (.A0(\efabless_subsystem.imem_wdata[0] ),
    .A1(\efabless_subsystem._003_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g197._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g197._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g197._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g2._1_  (.A0(\efabless_subsystem.imem_wdata[195] ),
    .A1(\efabless_subsystem._198_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g2._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[195] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g20._1_  (.A0(\efabless_subsystem.imem_wdata[177] ),
    .A1(\efabless_subsystem._180_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g20._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g20._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g20._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[177] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g21._1_  (.A0(\efabless_subsystem.imem_wdata[176] ),
    .A1(\efabless_subsystem._179_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g21._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g21._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g21._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[176] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g22._1_  (.A0(\efabless_subsystem.imem_wdata[175] ),
    .A1(\efabless_subsystem._178_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g22._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g22._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g22._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[175] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g23._1_  (.A0(\efabless_subsystem.imem_wdata[174] ),
    .A1(\efabless_subsystem._177_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g23._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g23._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g23._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[174] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g24._1_  (.A0(\efabless_subsystem.imem_wdata[173] ),
    .A1(\efabless_subsystem._176_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g24._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[173] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g25._1_  (.A0(\efabless_subsystem.imem_wdata[172] ),
    .A1(\efabless_subsystem._175_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g25._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[172] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g26._1_  (.A0(\efabless_subsystem.imem_wdata[171] ),
    .A1(\efabless_subsystem._174_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g26._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g26._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g26._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[171] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g27._1_  (.A0(\efabless_subsystem.imem_wdata[170] ),
    .A1(\efabless_subsystem._173_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g27._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g27._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g27._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[170] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g28._1_  (.A0(\efabless_subsystem.imem_wdata[169] ),
    .A1(\efabless_subsystem._172_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g28._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g28._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g28._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[169] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g29._1_  (.A0(\efabless_subsystem.imem_wdata[168] ),
    .A1(\efabless_subsystem._171_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g29._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g29._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g29._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[168] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g3._1_  (.A0(\efabless_subsystem.imem_wdata[194] ),
    .A1(\efabless_subsystem._197_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g3._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[194] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g30._1_  (.A0(\efabless_subsystem.imem_wdata[167] ),
    .A1(\efabless_subsystem._170_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g30._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g30._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g30._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[167] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g31._1_  (.A0(\efabless_subsystem.imem_wdata[166] ),
    .A1(\efabless_subsystem._169_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g31._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g31._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g31._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[166] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g32._1_  (.A0(\efabless_subsystem.imem_wdata[165] ),
    .A1(\efabless_subsystem._168_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g32._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[165] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g33._1_  (.A0(\efabless_subsystem.imem_wdata[164] ),
    .A1(\efabless_subsystem._167_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g33._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g33._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g33._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[164] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g34._1_  (.A0(\efabless_subsystem.imem_wdata[163] ),
    .A1(\efabless_subsystem._166_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g34._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g34._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g34._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[163] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g35._1_  (.A0(\efabless_subsystem.imem_wdata[162] ),
    .A1(\efabless_subsystem._165_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g35._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g35._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g35._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[162] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g36._1_  (.A0(\efabless_subsystem.imem_wdata[161] ),
    .A1(\efabless_subsystem._164_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g36._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g36._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g36._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[161] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g37._1_  (.A0(\efabless_subsystem.imem_wdata[160] ),
    .A1(\efabless_subsystem._163_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g37._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g37._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g37._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[160] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g38._1_  (.A0(\efabless_subsystem.imem_wdata[159] ),
    .A1(\efabless_subsystem._162_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g38._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g38._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g38._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[159] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g39._1_  (.A0(\efabless_subsystem.imem_wdata[158] ),
    .A1(\efabless_subsystem._161_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g39._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g39._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g39._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[158] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g4._1_  (.A0(\efabless_subsystem.imem_wdata[193] ),
    .A1(\efabless_subsystem._196_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g4._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[193] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g40._1_  (.A0(\efabless_subsystem.imem_wdata[157] ),
    .A1(\efabless_subsystem._160_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g40._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g40._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g40._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[157] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g41._1_  (.A0(\efabless_subsystem.imem_wdata[156] ),
    .A1(\efabless_subsystem._159_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g41._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g41._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g41._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[156] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g42._1_  (.A0(\efabless_subsystem.imem_wdata[155] ),
    .A1(\efabless_subsystem._158_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g42._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g42._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g42._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[155] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g43._1_  (.A0(\efabless_subsystem.imem_wdata[154] ),
    .A1(\efabless_subsystem._157_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g43._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g43._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g43._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[154] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g44._1_  (.A0(\efabless_subsystem.imem_wdata[153] ),
    .A1(\efabless_subsystem._156_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g44._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g44._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g44._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[153] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g45._1_  (.A0(\efabless_subsystem.imem_wdata[152] ),
    .A1(\efabless_subsystem._155_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g45._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g45._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g45._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[152] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g46._1_  (.A0(\efabless_subsystem.imem_wdata[151] ),
    .A1(\efabless_subsystem._154_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g46._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g46._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g46._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[151] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g47._1_  (.A0(\efabless_subsystem.imem_wdata[150] ),
    .A1(\efabless_subsystem._153_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g47._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g47._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g47._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[150] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g48._1_  (.A0(\efabless_subsystem.imem_wdata[149] ),
    .A1(\efabless_subsystem._152_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g48._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g48._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g48._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[149] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g49._1_  (.A0(\efabless_subsystem.imem_wdata[148] ),
    .A1(\efabless_subsystem._151_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g49._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g49._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g49._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[148] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g5._1_  (.A0(\efabless_subsystem.imem_wdata[192] ),
    .A1(\efabless_subsystem._195_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g5._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[192] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g50._1_  (.A0(\efabless_subsystem.imem_wdata[147] ),
    .A1(\efabless_subsystem._150_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g50._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g50._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g50._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[147] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g51._1_  (.A0(\efabless_subsystem.imem_wdata[146] ),
    .A1(\efabless_subsystem._149_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g51._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g51._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g51._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[146] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g52._1_  (.A0(\efabless_subsystem.imem_wdata[145] ),
    .A1(\efabless_subsystem._148_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g52._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g52._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g52._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[145] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g53._1_  (.A0(\efabless_subsystem.imem_wdata[144] ),
    .A1(\efabless_subsystem._147_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g53._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g53._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g53._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[144] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g54._1_  (.A0(\efabless_subsystem.imem_wdata[143] ),
    .A1(\efabless_subsystem._146_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g54._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g54._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g54._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[143] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g55._1_  (.A0(\efabless_subsystem.imem_wdata[142] ),
    .A1(\efabless_subsystem._145_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g55._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g55._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g55._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[142] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g56._1_  (.A0(\efabless_subsystem.imem_wdata[141] ),
    .A1(\efabless_subsystem._144_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g56._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g56._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g56._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[141] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g57._1_  (.A0(\efabless_subsystem.imem_wdata[140] ),
    .A1(\efabless_subsystem._143_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g57._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g57._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g57._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[140] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g58._1_  (.A0(\efabless_subsystem.imem_wdata[139] ),
    .A1(\efabless_subsystem._142_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g58._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g58._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g58._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[139] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g59._1_  (.A0(\efabless_subsystem.imem_wdata[138] ),
    .A1(\efabless_subsystem._141_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g59._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g59._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g59._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[138] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g6._1_  (.A0(\efabless_subsystem.imem_wdata[191] ),
    .A1(\efabless_subsystem._194_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g6._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[191] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g60._1_  (.A0(\efabless_subsystem.imem_wdata[137] ),
    .A1(\efabless_subsystem._140_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g60._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g60._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g60._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[137] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g61._1_  (.A0(\efabless_subsystem.imem_wdata[136] ),
    .A1(\efabless_subsystem._139_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g61._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g61._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g61._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[136] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g62._1_  (.A0(\efabless_subsystem.imem_wdata[135] ),
    .A1(\efabless_subsystem._138_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g62._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g62._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g62._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[135] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g63._1_  (.A0(\efabless_subsystem.imem_wdata[134] ),
    .A1(\efabless_subsystem._137_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g63._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g63._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g63._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[134] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g64._1_  (.A0(\efabless_subsystem.imem_wdata[133] ),
    .A1(\efabless_subsystem._136_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g64._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g64._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g64._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[133] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g65._1_  (.A0(\efabless_subsystem.imem_wdata[132] ),
    .A1(\efabless_subsystem._135_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g65._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g65._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g65._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[132] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g66._1_  (.A0(\efabless_subsystem.imem_wdata[131] ),
    .A1(\efabless_subsystem._134_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g66._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g66._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g66._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[131] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g67._1_  (.A0(\efabless_subsystem.imem_wdata[130] ),
    .A1(\efabless_subsystem._133_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g67._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g67._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g67._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[130] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g68._1_  (.A0(\efabless_subsystem.imem_wdata[129] ),
    .A1(\efabless_subsystem._132_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g68._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g68._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g68._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[129] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g69._1_  (.A0(\efabless_subsystem.imem_wdata[128] ),
    .A1(\efabless_subsystem._131_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g69._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g69._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g69._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[128] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g7._1_  (.A0(\efabless_subsystem.imem_wdata[190] ),
    .A1(\efabless_subsystem._193_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[190] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g70._1_  (.A0(\efabless_subsystem.imem_wdata[127] ),
    .A1(\efabless_subsystem._130_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g70._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g70._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g70._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[127] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g71._1_  (.A0(\efabless_subsystem.imem_wdata[126] ),
    .A1(\efabless_subsystem._129_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g71._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g71._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g71._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[126] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g72._1_  (.A0(\efabless_subsystem.imem_wdata[125] ),
    .A1(\efabless_subsystem._128_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g72._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g72._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g72._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[125] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g73._1_  (.A0(\efabless_subsystem.imem_wdata[124] ),
    .A1(\efabless_subsystem._127_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g73._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g73._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g73._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[124] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g74._1_  (.A0(\efabless_subsystem.imem_wdata[123] ),
    .A1(\efabless_subsystem._126_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g74._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g74._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g74._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[123] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g75._1_  (.A0(\efabless_subsystem.imem_wdata[122] ),
    .A1(\efabless_subsystem._125_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g75._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g75._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g75._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[122] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g76._1_  (.A0(\efabless_subsystem.imem_wdata[121] ),
    .A1(\efabless_subsystem._124_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g76._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g76._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g76._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[121] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g77._1_  (.A0(\efabless_subsystem.imem_wdata[120] ),
    .A1(\efabless_subsystem._123_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g77._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g77._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g77._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[120] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g78._1_  (.A0(\efabless_subsystem.imem_wdata[119] ),
    .A1(\efabless_subsystem._122_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g78._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g78._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g78._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[119] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g79._1_  (.A0(\efabless_subsystem.imem_wdata[118] ),
    .A1(\efabless_subsystem._121_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g79._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g79._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g79._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[118] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g8._1_  (.A0(\efabless_subsystem.imem_wdata[189] ),
    .A1(\efabless_subsystem._192_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[189] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g80._1_  (.A0(\efabless_subsystem.imem_wdata[117] ),
    .A1(\efabless_subsystem._120_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g80._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g80._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g80._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[117] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g81._1_  (.A0(\efabless_subsystem.imem_wdata[116] ),
    .A1(\efabless_subsystem._119_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g81._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g81._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g81._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[116] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g82._1_  (.A0(\efabless_subsystem.imem_wdata[115] ),
    .A1(\efabless_subsystem._118_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g82._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g82._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g82._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[115] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g83._1_  (.A0(\efabless_subsystem.imem_wdata[114] ),
    .A1(\efabless_subsystem._117_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g83._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g83._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g83._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[114] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g84._1_  (.A0(\efabless_subsystem.imem_wdata[113] ),
    .A1(\efabless_subsystem._116_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g84._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g84._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g84._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[113] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g85._1_  (.A0(\efabless_subsystem.imem_wdata[112] ),
    .A1(\efabless_subsystem._115_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g85._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g85._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g85._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[112] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g86._1_  (.A0(\efabless_subsystem.imem_wdata[111] ),
    .A1(\efabless_subsystem._114_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g86._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g86._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g86._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[111] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g87._1_  (.A0(\efabless_subsystem.imem_wdata[110] ),
    .A1(\efabless_subsystem._113_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g87._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g87._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g87._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[110] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g88._1_  (.A0(\efabless_subsystem.imem_wdata[109] ),
    .A1(\efabless_subsystem._112_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g88._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g88._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g88._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[109] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g89._1_  (.A0(\efabless_subsystem.imem_wdata[108] ),
    .A1(\efabless_subsystem._111_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g89._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g89._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g89._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[108] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g9._1_  (.A0(\efabless_subsystem.imem_wdata[188] ),
    .A1(\efabless_subsystem._191_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[188] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g90._1_  (.A0(\efabless_subsystem.imem_wdata[107] ),
    .A1(\efabless_subsystem._110_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g90._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g90._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g90._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[107] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g91._1_  (.A0(\efabless_subsystem.imem_wdata[106] ),
    .A1(\efabless_subsystem._109_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g91._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g91._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g91._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[106] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g92._1_  (.A0(\efabless_subsystem.imem_wdata[105] ),
    .A1(\efabless_subsystem._108_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g92._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g92._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g92._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[105] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g93._1_  (.A0(\efabless_subsystem.imem_wdata[104] ),
    .A1(\efabless_subsystem._107_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g93._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g93._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g93._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[104] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g94._1_  (.A0(\efabless_subsystem.imem_wdata[103] ),
    .A1(\efabless_subsystem._106_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g94._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g94._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g94._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[103] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g95._1_  (.A0(\efabless_subsystem.imem_wdata[102] ),
    .A1(\efabless_subsystem._105_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g95._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g95._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g95._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[102] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g96._1_  (.A0(\efabless_subsystem.imem_wdata[101] ),
    .A1(\efabless_subsystem._104_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g96._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g96._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g96._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[101] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g97._1_  (.A0(\efabless_subsystem.imem_wdata[100] ),
    .A1(\efabless_subsystem._103_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g97._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g97._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g97._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[100] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g98._1_  (.A0(\efabless_subsystem.imem_wdata[99] ),
    .A1(\efabless_subsystem._102_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g98._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g98._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g98._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[99] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_82_26.g99._1_  (.A0(\efabless_subsystem.imem_wdata[98] ),
    .A1(\efabless_subsystem._101_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_82_26.g99._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_82_26.g99._2_  (.A(\efabless_subsystem.input_memory_i.mux_82_26.g99._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wdata[98] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g1._1_  (.A0(\efabless_subsystem.imem_wmask[192] ),
    .A1(\efabless_subsystem.input_memory_i._037_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[24] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g10._1_  (.A0(\efabless_subsystem.imem_wmask[120] ),
    .A1(\efabless_subsystem.input_memory_i._028_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[15] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g11._1_  (.A0(\efabless_subsystem.imem_wmask[112] ),
    .A1(\efabless_subsystem.input_memory_i._027_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[14] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g12._1_  (.A0(\efabless_subsystem.imem_wmask[104] ),
    .A1(\efabless_subsystem.input_memory_i._026_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[13] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g13._1_  (.A0(\efabless_subsystem.imem_wmask[96] ),
    .A1(\efabless_subsystem.input_memory_i._025_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g13._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[12] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g14._1_  (.A0(\efabless_subsystem.imem_wmask[88] ),
    .A1(\efabless_subsystem.input_memory_i._024_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g14._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[11] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g15._1_  (.A0(\efabless_subsystem.imem_wmask[80] ),
    .A1(\efabless_subsystem.input_memory_i._023_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g15._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[10] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g16._1_  (.A0(\efabless_subsystem.imem_wmask[72] ),
    .A1(\efabless_subsystem.input_memory_i._022_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g16._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[9] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g17._1_  (.A0(\efabless_subsystem.imem_wmask[64] ),
    .A1(\efabless_subsystem.input_memory_i._021_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g17._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g17._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g17._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[8] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g18._1_  (.A0(\efabless_subsystem.imem_wmask[56] ),
    .A1(\efabless_subsystem.input_memory_i._020_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g18._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g18._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g18._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[7] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g19._1_  (.A0(\efabless_subsystem.imem_wmask[48] ),
    .A1(\efabless_subsystem.input_memory_i._019_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g19._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g19._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g19._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[6] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g2._1_  (.A0(\efabless_subsystem.imem_wmask[184] ),
    .A1(\efabless_subsystem.input_memory_i._036_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g2._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[23] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g20._1_  (.A0(\efabless_subsystem.imem_wmask[40] ),
    .A1(\efabless_subsystem.input_memory_i._018_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g20._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g20._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g20._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[5] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g21._1_  (.A0(\efabless_subsystem.imem_wmask[32] ),
    .A1(\efabless_subsystem.input_memory_i._017_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g21._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g21._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g21._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g22._1_  (.A0(\efabless_subsystem.imem_wmask[24] ),
    .A1(\efabless_subsystem.input_memory_i._016_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g22._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g22._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g22._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g23._1_  (.A0(\efabless_subsystem.imem_wmask[16] ),
    .A1(\efabless_subsystem.input_memory_i._015_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g23._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g23._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g23._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g24._1_  (.A0(\efabless_subsystem.imem_wmask[8] ),
    .A1(\efabless_subsystem.input_memory_i._014_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g24._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g25._1_  (.A0(\efabless_subsystem.imem_wmask[0] ),
    .A1(\efabless_subsystem.input_memory_i._013_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g25._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g25._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g25._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g3._1_  (.A0(\efabless_subsystem.imem_wmask[176] ),
    .A1(\efabless_subsystem.input_memory_i._035_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g3._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[22] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g4._1_  (.A0(\efabless_subsystem.imem_wmask[168] ),
    .A1(\efabless_subsystem.input_memory_i._034_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g4._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[21] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g5._1_  (.A0(\efabless_subsystem.imem_wmask[160] ),
    .A1(\efabless_subsystem.input_memory_i._033_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g5._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[20] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g6._1_  (.A0(\efabless_subsystem.imem_wmask[152] ),
    .A1(\efabless_subsystem.input_memory_i._032_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g6._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[19] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g7._1_  (.A0(\efabless_subsystem.imem_wmask[144] ),
    .A1(\efabless_subsystem.input_memory_i._031_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[18] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g8._1_  (.A0(\efabless_subsystem.imem_wmask[136] ),
    .A1(\efabless_subsystem.input_memory_i._030_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[17] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_83_26.g9._1_  (.A0(\efabless_subsystem.imem_wmask[128] ),
    .A1(\efabless_subsystem.input_memory_i._029_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_83_26.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_83_26.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_83_26.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wmask[16] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_84_26.g10._1_  (.A0(\efabless_subsystem.imem_address[2] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_84_26.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_84_26.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_84_26.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_addr[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_84_26.g11._1_  (.A0(\efabless_subsystem.imem_address[1] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_84_26.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_84_26.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_84_26.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_addr[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_84_26.g12._1_  (.A0(\efabless_subsystem.imem_address[0] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_84_26.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_84_26.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_84_26.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_addr[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_84_26.g7._1_  (.A0(\efabless_subsystem.imem_address[5] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_84_26.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_84_26.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_84_26.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_addr[5] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_84_26.g8._1_  (.A0(\efabless_subsystem.imem_address[4] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_84_26.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_84_26.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_84_26.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_addr[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_84_26.g9._1_  (.A0(\efabless_subsystem.imem_address[3] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_84_26.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_84_26.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_84_26.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_addr[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_85_26.g1._1_  (.A0(\efabless_subsystem.imem_wren ),
    .A1(\efabless_subsystem.input_memory_i.mux_85_26.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_85_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_85_26.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_85_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.memory_wren ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.input_memory_i.mux_fifo_state_103_19.g1._0_  (.A1(\efabless_subsystem.input_memory_i._038_ ),
    .A2(\efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[1] ),
    .B1(\efabless_subsystem.input_memory_i._083_ ),
    .B2(\efabless_subsystem.input_memory_i.ctl_fifo_state_103_19.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.fifo_state_reg[0].d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[12] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[3] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[2] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[1] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[0] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[11] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[10] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[9] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[8] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[7] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[6] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[5] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9._1_  (.A0(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_rdptr_init[4] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g1._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[12] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[12] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g10._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[3] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g11._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[2] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g12._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[1] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g13._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[0] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g13._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g2._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[11] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g2._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g3._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[10] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g3._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g4._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[9] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g4._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g5._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[8] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g5._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g6._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[7] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g6._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g7._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[6] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g8._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[5] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g9._1_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .A1(\efabless_subsystem.input_memory_i.add_149_37.Z[4] ),
    .S(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_read_ptr_d_148_22.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[12] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[3] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[2] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[1] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[0] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[11] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[10] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[9] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[8] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[7] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[6] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[5] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9._1_  (.A0(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_imem_fifo_wrptr_init[4] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g1._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[12] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[12] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g1._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g10._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[3] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g10._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g11._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[2] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g11._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g12._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[1] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g12._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g13._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[0] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g13._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g2._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[11] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g2._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g3._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[10] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g3._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g4._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[9] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g4._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g5._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[8] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g5._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g6._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[7] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g6._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g7._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[6] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g7._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g8._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[5] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g8._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g9._1_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .A1(\efabless_subsystem.input_memory_i.add_144_39.Z[4] ),
    .S(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g9._2_  (.A(\efabless_subsystem.input_memory_i.mux_write_ptr_d_143_33.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9.data0 ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._00_ ),
    .B(\efabless_subsystem.input_memory_i._084_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g13.z ),
    .S(\efabless_subsystem.input_memory_i._039_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._085_ ),
    .S(\efabless_subsystem.input_memory_i._086_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[0] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._00_ ),
    .B(\efabless_subsystem.input_memory_i._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g3.z ),
    .S(\efabless_subsystem.input_memory_i._040_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._088_ ),
    .S(\efabless_subsystem.input_memory_i._089_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[10] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._00_ ),
    .B(\efabless_subsystem.input_memory_i._090_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g2.z ),
    .S(\efabless_subsystem.input_memory_i._041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._091_ ),
    .S(\efabless_subsystem.input_memory_i._092_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[11] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._00_ ),
    .B(\efabless_subsystem.input_memory_i._093_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[12] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g1.z ),
    .S(\efabless_subsystem.input_memory_i._042_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._094_ ),
    .S(\efabless_subsystem.input_memory_i._095_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[12] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._00_ ),
    .B(\efabless_subsystem.input_memory_i._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g12.z ),
    .S(\efabless_subsystem.input_memory_i._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._097_ ),
    .S(\efabless_subsystem.input_memory_i._098_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[1] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._00_ ),
    .B(\efabless_subsystem.input_memory_i._099_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g11.z ),
    .S(\efabless_subsystem.input_memory_i._044_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._100_ ),
    .S(\efabless_subsystem.input_memory_i._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[2] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._00_ ),
    .B(\efabless_subsystem.input_memory_i._102_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g10.z ),
    .S(\efabless_subsystem.input_memory_i._045_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._103_ ),
    .S(\efabless_subsystem.input_memory_i._104_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[3] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._00_ ),
    .B(\efabless_subsystem.input_memory_i._105_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g9.z ),
    .S(\efabless_subsystem.input_memory_i._046_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._106_ ),
    .S(\efabless_subsystem.input_memory_i._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[4] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._00_ ),
    .B(\efabless_subsystem.input_memory_i._108_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g8.z ),
    .S(\efabless_subsystem.input_memory_i._047_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._109_ ),
    .S(\efabless_subsystem.input_memory_i._110_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[5] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._00_ ),
    .B(\efabless_subsystem.input_memory_i._111_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g7.z ),
    .S(\efabless_subsystem.input_memory_i._048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._112_ ),
    .S(\efabless_subsystem.input_memory_i._113_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[6] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._00_ ),
    .B(\efabless_subsystem.input_memory_i._114_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g6.z ),
    .S(\efabless_subsystem.input_memory_i._049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._115_ ),
    .S(\efabless_subsystem.input_memory_i._116_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[7] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._00_ ),
    .B(\efabless_subsystem.input_memory_i._117_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g5.z ),
    .S(\efabless_subsystem.input_memory_i._050_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._118_ ),
    .S(\efabless_subsystem.input_memory_i._119_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[8] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._08_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._00_ ),
    .B(\efabless_subsystem.input_memory_i._120_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._09_  (.A0(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .A1(\efabless_subsystem.input_memory_i.mux_read_ptr_d_135_9.g4.z ),
    .S(\efabless_subsystem.input_memory_i._051_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._10_  (.A0(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._121_ ),
    .S(\efabless_subsystem.input_memory_i._122_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._11_  (.A(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._02_ ),
    .D(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_149_37.A[9] ),
    .Q_N(\efabless_subsystem.input_memory_i.read_ptr_q_reg[9]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._00_ ),
    .B(\efabless_subsystem.input_memory_i._123_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g13.z ),
    .S(\efabless_subsystem.input_memory_i._052_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._124_ ),
    .S(\efabless_subsystem.input_memory_i._125_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[0] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._00_ ),
    .B(\efabless_subsystem.input_memory_i._126_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g3.z ),
    .S(\efabless_subsystem.input_memory_i._053_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._127_ ),
    .S(\efabless_subsystem.input_memory_i._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[10] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[10]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._00_ ),
    .B(\efabless_subsystem.input_memory_i._129_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g2.z ),
    .S(\efabless_subsystem.input_memory_i._054_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._130_ ),
    .S(\efabless_subsystem.input_memory_i._131_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[11] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[11]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._00_ ),
    .B(\efabless_subsystem.input_memory_i._132_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[12] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g1.z ),
    .S(\efabless_subsystem.input_memory_i._055_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._133_ ),
    .S(\efabless_subsystem.input_memory_i._134_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[12] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[12]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._00_ ),
    .B(\efabless_subsystem.input_memory_i._135_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g12.z ),
    .S(\efabless_subsystem.input_memory_i._056_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._136_ ),
    .S(\efabless_subsystem.input_memory_i._137_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[1] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._00_ ),
    .B(\efabless_subsystem.input_memory_i._138_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g11.z ),
    .S(\efabless_subsystem.input_memory_i._057_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._139_ ),
    .S(\efabless_subsystem.input_memory_i._140_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[2] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._00_ ),
    .B(\efabless_subsystem.input_memory_i._141_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g10.z ),
    .S(\efabless_subsystem.input_memory_i._058_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._142_ ),
    .S(\efabless_subsystem.input_memory_i._143_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[3] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._00_ ),
    .B(\efabless_subsystem.input_memory_i._144_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g9.z ),
    .S(\efabless_subsystem.input_memory_i._059_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._145_ ),
    .S(\efabless_subsystem.input_memory_i._146_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[4] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._00_ ),
    .B(\efabless_subsystem.input_memory_i._147_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g8.z ),
    .S(\efabless_subsystem.input_memory_i._060_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._148_ ),
    .S(\efabless_subsystem.input_memory_i._149_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[5] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._00_ ),
    .B(\efabless_subsystem.input_memory_i._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g7.z ),
    .S(\efabless_subsystem.input_memory_i._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._151_ ),
    .S(\efabless_subsystem.input_memory_i._152_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[6] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._00_ ),
    .B(\efabless_subsystem.input_memory_i._153_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g6.z ),
    .S(\efabless_subsystem.input_memory_i._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._154_ ),
    .S(\efabless_subsystem.input_memory_i._155_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[7] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._00_ ),
    .B(\efabless_subsystem.input_memory_i._156_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g5.z ),
    .S(\efabless_subsystem.input_memory_i._063_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._157_ ),
    .S(\efabless_subsystem.input_memory_i._158_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[8] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._07_  (.A(\efabless_subsystem.input_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._08_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._00_ ),
    .B(\efabless_subsystem.input_memory_i._159_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._09_  (.A0(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .A1(\efabless_subsystem.input_memory_i.mux_write_ptr_d_135_9.g4.z ),
    .S(\efabless_subsystem.input_memory_i._064_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._10_  (.A0(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._04_ ),
    .A1(\efabless_subsystem.input_memory_i._160_ ),
    .S(\efabless_subsystem.input_memory_i._161_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._11_  (.A(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._13_  (.CLK_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._02_ ),
    .D(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._03_ ),
    .RESET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._00_ ),
    .SET_B(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.input_memory_i.add_144_39.A[9] ),
    .Q_N(\efabless_subsystem.input_memory_i.write_ptr_q_reg[9]._06_ ));
 sky130_fd_sc_hd__nor4_2 \efabless_subsystem.mmap_interconnect_i._0314_  (.A(\efabless_subsystem.cpu_address[22] ),
    .B(\efabless_subsystem.cpu_address[23] ),
    .C(\efabless_subsystem.cpu_address[21] ),
    .D(\efabless_subsystem.cpu_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_105_36.ctl ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.mmap_interconnect_i._0315_  (.A_N(\efabless_subsystem.cpu_address[2] ),
    .B(\efabless_subsystem.cpu_address[3] ),
    .C(\efabless_subsystem.cpu_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i._0000_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i._0316_  (.A(\efabless_subsystem.mmap_interconnect_i._0000_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.ctl ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.mmap_interconnect_i._0317_  (.A_N(\efabless_subsystem.cpu_address[3] ),
    .B(\efabless_subsystem.cpu_address[4] ),
    .C(\efabless_subsystem.cpu_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i._0001_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i._0318_  (.A(\efabless_subsystem.mmap_interconnect_i._0001_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.ctl ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.mmap_interconnect_i._0319_  (.A(\efabless_subsystem.cpu_address[2] ),
    .B(\efabless_subsystem.cpu_address[3] ),
    .C_N(\efabless_subsystem.cpu_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.ctl ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.mmap_interconnect_i._0320_  (.A_N(\efabless_subsystem.cpu_address[4] ),
    .B(\efabless_subsystem.cpu_address[3] ),
    .C(\efabless_subsystem.cpu_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i._0002_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i._0321_  (.A(\efabless_subsystem.mmap_interconnect_i._0002_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.ctl ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.mmap_interconnect_i._0322_  (.A(\efabless_subsystem.cpu_address[2] ),
    .B(\efabless_subsystem.cpu_address[4] ),
    .C_N(\efabless_subsystem.cpu_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.ctl ));
 sky130_fd_sc_hd__nor3b_2 \efabless_subsystem.mmap_interconnect_i._0323_  (.A(\efabless_subsystem.cpu_address[3] ),
    .B(\efabless_subsystem.cpu_address[4] ),
    .C_N(\efabless_subsystem.cpu_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.ctl ));
 sky130_fd_sc_hd__nor3_2 \efabless_subsystem.mmap_interconnect_i._0324_  (.A(\efabless_subsystem.cpu_address[2] ),
    .B(\efabless_subsystem.cpu_address[3] ),
    .C(\efabless_subsystem.cpu_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.ctl ));
 sky130_fd_sc_hd__nor4b_2 \efabless_subsystem.mmap_interconnect_i._0325_  (.A(\efabless_subsystem.cpu_address[22] ),
    .B(\efabless_subsystem.cpu_address[23] ),
    .C(\efabless_subsystem.cpu_address[21] ),
    .D_N(\efabless_subsystem.cpu_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_106_36.ctl ));
 sky130_fd_sc_hd__nor4b_2 \efabless_subsystem.mmap_interconnect_i._0326_  (.A(\efabless_subsystem.cpu_address[22] ),
    .B(\efabless_subsystem.cpu_address[23] ),
    .C(\efabless_subsystem.cpu_address[20] ),
    .D_N(\efabless_subsystem.cpu_address[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.mmap_interconnect_i.mux_107_36.ctl ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0329_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0004_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0330_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0005_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0331_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0006_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0334_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0009_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0335_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0010_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0364_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0039_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0372_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0380_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0055_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0388_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0063_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0396_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0071_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0404_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0412_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0087_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0420_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0428_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0103_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0436_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0111_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0444_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0119_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0452_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0127_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0460_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0135_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0468_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0143_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0476_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0151_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0484_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0159_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0492_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0167_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0500_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0175_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0508_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0183_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0516_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0191_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0524_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0199_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0556_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0231_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0564_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0239_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0572_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0247_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.mmap_interconnect_i._0580_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.mmap_interconnect_i._0255_ ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0649_  (.A(\efabless_subsystem.cpu_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0650_  (.A(\efabless_subsystem.cpu_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0651_  (.A(\efabless_subsystem.cpu_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0652_  (.A(\efabless_subsystem.cpu_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0653_  (.A(\efabless_subsystem.cpu_address[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0654_  (.A(\efabless_subsystem.cpu_address[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0655_  (.A(\efabless_subsystem.cpu_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0656_  (.A(\efabless_subsystem.cpu_address[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0657_  (.A(\efabless_subsystem.cpu_address[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0658_  (.A(\efabless_subsystem.cpu_address[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0659_  (.A(\efabless_subsystem.cpu_address[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0660_  (.A(\efabless_subsystem.cpu_address[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0661_  (.A(\efabless_subsystem.cpu_address[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0662_  (.A(\efabless_subsystem.cpu_address[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0663_  (.A(\efabless_subsystem.cpu_address[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0664_  (.A(\efabless_subsystem.cpu_address[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0665_  (.A(\efabless_subsystem.cpu_address[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0666_  (.A(\efabless_subsystem.cpu_address[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0667_  (.A(\efabless_subsystem.cpu_address[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0668_  (.A(\efabless_subsystem.cpu_address[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0669_  (.A(\efabless_subsystem.cpu_address[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0670_  (.A(\efabless_subsystem.cpu_address[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_address[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0679_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0680_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0681_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0682_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0683_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0684_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0685_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0686_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0687_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0688_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0689_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0690_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0691_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0692_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0693_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0694_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0695_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0696_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0697_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0698_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0699_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0700_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0701_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0702_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0703_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0704_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0705_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0706_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0707_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0708_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0709_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[30] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0710_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_data_in[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0711_  (.A(\efabless_subsystem.cpu_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0712_  (.A(\efabless_subsystem.cpu_wmask[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0713_  (.A(\efabless_subsystem.cpu_wmask[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0714_  (.A(\efabless_subsystem.cpu_wmask[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0715_  (.A(\efabless_subsystem.cpu_wmask[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0716_  (.A(\efabless_subsystem.cpu_wmask[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0717_  (.A(\efabless_subsystem.cpu_wmask[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0718_  (.A(\efabless_subsystem.cpu_wmask[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0719_  (.A(\efabless_subsystem.cpu_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0720_  (.A(\efabless_subsystem.cpu_wmask[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0721_  (.A(\efabless_subsystem.cpu_wmask[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0722_  (.A(\efabless_subsystem.cpu_wmask[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0723_  (.A(\efabless_subsystem.cpu_wmask[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0724_  (.A(\efabless_subsystem.cpu_wmask[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0725_  (.A(\efabless_subsystem.cpu_wmask[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0726_  (.A(\efabless_subsystem.cpu_wmask[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0727_  (.A(\efabless_subsystem.cpu_wmask[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0728_  (.A(\efabless_subsystem.cpu_wmask[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0729_  (.A(\efabless_subsystem.cpu_wmask[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0730_  (.A(\efabless_subsystem.cpu_wmask[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0731_  (.A(\efabless_subsystem.cpu_wmask[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0732_  (.A(\efabless_subsystem.cpu_wmask[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0733_  (.A(\efabless_subsystem.cpu_wmask[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0734_  (.A(\efabless_subsystem.cpu_wmask[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0735_  (.A(\efabless_subsystem.cpu_wmask[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0736_  (.A(\efabless_subsystem.cpu_wmask[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0737_  (.A(\efabless_subsystem.cpu_wmask[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0738_  (.A(\efabless_subsystem.cpu_wmask[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0739_  (.A(\efabless_subsystem.cpu_wmask[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0740_  (.A(\efabless_subsystem.cpu_wmask[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0741_  (.A(\efabless_subsystem.cpu_wmask[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[30] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0742_  (.A(\efabless_subsystem.cpu_wmask[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wmask[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0743_  (.A(\efabless_subsystem.cpu_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_address[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0744_  (.A(\efabless_subsystem.cpu_address[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_address[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0745_  (.A(\efabless_subsystem.cpu_address[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_address[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0746_  (.A(\efabless_subsystem.cpu_address[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_address[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0747_  (.A(\efabless_subsystem.cpu_address[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_address[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0748_  (.A(\efabless_subsystem.cpu_address[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_address[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0770_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0771_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0772_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0773_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0774_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0775_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0776_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0777_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0778_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0779_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0780_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0781_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0782_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0783_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0784_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0785_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0786_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0787_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0788_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0789_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0790_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0791_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0792_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0793_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0794_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0795_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0796_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0797_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0798_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0799_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0800_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[30] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0801_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0802_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[32] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0803_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[33] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0804_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[34] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0805_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[35] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0806_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[36] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0807_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[37] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0808_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[38] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0809_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[39] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0810_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[40] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0811_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[41] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0812_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[42] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0813_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[43] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0814_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[44] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0815_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[45] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0816_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[46] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0817_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[47] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0818_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[48] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0819_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[49] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0820_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[50] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0821_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[51] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0822_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[52] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0823_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[53] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0824_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[54] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0825_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[55] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0826_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[56] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0827_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[57] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0828_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[58] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0829_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[59] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0830_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[60] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0831_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[61] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0832_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[62] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0833_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[63] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0834_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[64] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0835_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[65] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0836_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[66] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0837_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[67] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0838_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[68] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0839_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[69] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0840_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[70] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0841_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[71] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0842_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[72] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0843_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[73] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0844_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[74] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0845_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[75] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0846_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[76] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0847_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[77] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0848_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[78] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0849_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[79] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0850_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[80] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0851_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[81] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0852_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[82] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0853_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[83] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0854_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[84] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0855_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[85] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0856_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[86] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0857_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[87] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0858_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[88] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0859_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[89] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0860_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[90] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0861_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[91] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0862_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[92] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0863_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[93] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0864_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[94] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0865_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[95] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0866_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[96] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0867_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[97] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0868_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[98] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0869_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[99] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0870_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[100] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0871_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[101] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0872_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[102] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0873_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[103] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0874_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[104] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0875_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[105] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0876_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[106] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0877_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[107] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0878_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[108] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0879_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[109] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0880_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[110] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0881_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[111] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0882_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[112] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0883_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[113] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0884_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[114] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0885_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[115] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0886_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[116] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0887_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[117] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0888_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[118] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0889_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[119] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0890_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[120] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0891_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[121] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0892_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[122] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0893_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[123] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0894_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[124] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0895_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[125] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0896_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[126] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0897_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[127] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0898_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[128] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0899_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[129] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0900_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[130] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0901_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[131] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0902_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[132] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0903_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[133] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0904_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[134] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0905_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[135] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0906_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[136] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0907_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[137] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0908_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[138] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0909_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[139] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0910_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[140] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0911_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[141] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0912_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[142] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0913_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[143] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0914_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[144] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0915_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[145] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0916_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[146] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0917_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[147] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0918_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[148] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0919_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[149] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0920_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[150] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0921_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[151] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0922_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[152] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0923_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[153] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0924_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[154] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0925_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[155] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0926_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[156] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0927_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[157] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0928_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[158] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0929_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[159] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0930_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[160] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0931_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[161] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0932_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[162] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0933_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[163] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0934_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[164] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0935_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[165] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0936_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[166] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0937_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[167] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0938_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[168] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0939_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[169] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0940_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[170] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0941_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[171] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0942_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[172] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0943_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[173] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0944_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[174] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0945_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[175] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0946_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[176] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0947_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[177] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0948_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[178] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0949_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[179] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0950_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[180] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0951_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[181] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0952_  (.A(\efabless_subsystem.cpu_wdata[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[182] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0953_  (.A(\efabless_subsystem.cpu_wdata[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[183] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0954_  (.A(\efabless_subsystem.cpu_wdata[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[184] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0955_  (.A(\efabless_subsystem.cpu_wdata[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[185] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0956_  (.A(\efabless_subsystem.cpu_wdata[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[186] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0957_  (.A(\efabless_subsystem.cpu_wdata[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[187] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0958_  (.A(\efabless_subsystem.cpu_wdata[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[188] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0959_  (.A(\efabless_subsystem.cpu_wdata[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[189] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0960_  (.A(\efabless_subsystem.cpu_wdata[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[190] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0961_  (.A(\efabless_subsystem.cpu_wdata[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[191] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0962_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[192] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0963_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[193] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0964_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[194] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0965_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[195] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._0966_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wdata[196] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1045_  (.A(\efabless_subsystem.cpu_address[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1046_  (.A(\efabless_subsystem.cpu_address[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1047_  (.A(\efabless_subsystem.cpu_address[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1048_  (.A(\efabless_subsystem.cpu_address[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1049_  (.A(\efabless_subsystem.cpu_address[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1075_  (.A(\efabless_subsystem.cpu_wdata[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1076_  (.A(\efabless_subsystem.cpu_wdata[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1077_  (.A(\efabless_subsystem.cpu_wdata[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1078_  (.A(\efabless_subsystem.cpu_wdata[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1079_  (.A(\efabless_subsystem.cpu_wdata[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1080_  (.A(\efabless_subsystem.cpu_wdata[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1081_  (.A(\efabless_subsystem.cpu_wdata[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1082_  (.A(\efabless_subsystem.cpu_wdata[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1083_  (.A(\efabless_subsystem.cpu_wdata[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1084_  (.A(\efabless_subsystem.cpu_wdata[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1085_  (.A(\efabless_subsystem.cpu_wdata[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1086_  (.A(\efabless_subsystem.cpu_wdata[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1087_  (.A(\efabless_subsystem.cpu_wdata[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1088_  (.A(\efabless_subsystem.cpu_wdata[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1089_  (.A(\efabless_subsystem.cpu_wdata[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1090_  (.A(\efabless_subsystem.cpu_wdata[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1091_  (.A(\efabless_subsystem.cpu_wdata[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1092_  (.A(\efabless_subsystem.cpu_wdata[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1093_  (.A(\efabless_subsystem.cpu_wdata[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1094_  (.A(\efabless_subsystem.cpu_wdata[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1095_  (.A(\efabless_subsystem.cpu_wdata[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1096_  (.A(\efabless_subsystem.cpu_wdata[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1097_  (.A(\efabless_subsystem.cpu_wmask[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1105_  (.A(\efabless_subsystem.cpu_wmask[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.mmap_interconnect_i._1113_  (.A(\efabless_subsystem.cpu_wmask[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[16] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_105_36.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0004_ ),
    .A1(\efabless_subsystem.cpu_wren ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_105_36.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_105_36.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_105_36.g1._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_105_36.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cfg_wren ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_106_36.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0005_ ),
    .A1(\efabless_subsystem.cpu_wren ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_106_36.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_106_36.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_106_36.g1._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_106_36.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wren ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_107_36.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0006_ ),
    .A1(\efabless_subsystem.cpu_wren ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_107_36.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_107_36.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_107_36.g1._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_107_36.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_107_36.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_111_36.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0009_ ),
    .A1(\efabless_subsystem.cpu_rden ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_106_36.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_111_36.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_111_36.g1._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_111_36.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_rden ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_112_36.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0010_ ),
    .A1(\efabless_subsystem.cpu_rden ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_107_36.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_112_36.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_112_36.g1._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_112_36.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_112_36.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0055_ ),
    .A1(\efabless_subsystem.cpu_wmask[16] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g16._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[48] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g24._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0047_ ),
    .A1(\efabless_subsystem.cpu_wmask[8] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g24._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[40] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0039_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[32] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0063_ ),
    .A1(\efabless_subsystem.cpu_wmask[24] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g8._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_11.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[56] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0087_ ),
    .A1(\efabless_subsystem.cpu_wmask[16] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g16._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[80] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g24._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0079_ ),
    .A1(\efabless_subsystem.cpu_wmask[8] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g24._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[72] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0071_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[64] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0095_ ),
    .A1(\efabless_subsystem.cpu_wmask[24] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g8._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_12.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[88] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0119_ ),
    .A1(\efabless_subsystem.cpu_wmask[16] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g16._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[112] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g24._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0111_ ),
    .A1(\efabless_subsystem.cpu_wmask[8] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g24._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[104] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0103_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[96] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0127_ ),
    .A1(\efabless_subsystem.cpu_wmask[24] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g8._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_13.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[120] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0151_ ),
    .A1(\efabless_subsystem.cpu_wmask[16] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g16._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[144] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g24._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0143_ ),
    .A1(\efabless_subsystem.cpu_wmask[8] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g24._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[136] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0135_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[128] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0159_ ),
    .A1(\efabless_subsystem.cpu_wmask[24] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g8._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_14.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[152] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0183_ ),
    .A1(\efabless_subsystem.cpu_wmask[16] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g16._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[176] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g24._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0175_ ),
    .A1(\efabless_subsystem.cpu_wmask[8] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g24._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[168] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0167_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[160] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0191_ ),
    .A1(\efabless_subsystem.cpu_wmask[24] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g8._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_15.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[184] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0199_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_16.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[192] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0247_ ),
    .A1(\efabless_subsystem.cpu_wmask[16] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g16._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[16] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g24._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0239_ ),
    .A1(\efabless_subsystem.cpu_wmask[8] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g24._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g24._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g24._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[8] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g32._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0231_ ),
    .A1(\efabless_subsystem.cpu_wmask[0] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g32._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g32._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g32._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i._0255_ ),
    .A1(\efabless_subsystem.cpu_wmask[24] ),
    .S(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g8._2_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_imem_wmask_expanded_181_35.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.imem_wmask[24] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mux_276_38.g1._1_  (.A0(\efabless_subsystem.compute_core_i.i_array_shftsgn_valid ),
    .A1(\efabless_subsystem.mux_276_38.g1.data1 ),
    .S(\efabless_subsystem.compute_core_i.i_stat_cfg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mux_276_38.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mux_276_38.g1._2_  (.A(\efabless_subsystem.mux_276_38.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.i_fmap_valid ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.mux_277_38.g1._1_  (.A0(\efabless_subsystem.mux_276_38.g1.data1 ),
    .A1(\efabless_subsystem.compute_core_i.i_array_shftsgn_valid ),
    .S(\efabless_subsystem.compute_core_i.i_stat_cfg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.mux_277_38.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.mux_277_38.g1._2_  (.A(\efabless_subsystem.mux_277_38.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.compute_core_i.i_weight_valid ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i._098_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i._099_  (.A(\efabless_subsystem.mmap_interconnect_i.mux_112_36.g1.z ),
    .B(\efabless_subsystem.reduction_memory_i.memory_wren ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.n_160 ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i._100_  (.A(\efabless_subsystem.reduction_memory_i.memory_wren ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.n_161 ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i._101_  (.A(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i._000_ ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.reduction_memory_i._102_  (.A(\efabless_subsystem.reduction_memory_i.g18.Z[4] ),
    .B(\efabless_subsystem.reduction_memory_i.g18.Z[2] ),
    .C(\efabless_subsystem.reduction_memory_i.g18.Z[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._001_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.reduction_memory_i._103_  (.A(\efabless_subsystem.reduction_memory_i.g18.Z[6] ),
    .B(\efabless_subsystem.reduction_memory_i.g18.Z[5] ),
    .C(\efabless_subsystem.reduction_memory_i.g18.Z[0] ),
    .D(\efabless_subsystem.reduction_memory_i.g18.Z[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._002_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.reduction_memory_i._104_  (.A(\efabless_subsystem.reduction_memory_i.g18.Z[7] ),
    .B(\efabless_subsystem.reduction_memory_i.g18.Z[8] ),
    .C(\efabless_subsystem.reduction_memory_i._001_ ),
    .D(\efabless_subsystem.reduction_memory_i._002_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._003_ ));
 sky130_fd_sc_hd__o21ai_2 \efabless_subsystem.reduction_memory_i._105_  (.A1(\efabless_subsystem.reduction_memory_i._000_ ),
    .A2(\efabless_subsystem.compute_controller_i.o_red_params_pop ),
    .B1(\efabless_subsystem.reduction_memory_i._003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.n_162 ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.reduction_memory_i._106_  (.A(\efabless_subsystem.compute_controller_i.o_red_params_pop ),
    .B(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._004_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i._107_  (.A0(\efabless_subsystem.reduction_memory_i._004_ ),
    .A1(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[1] ),
    .S(\efabless_subsystem.reduction_memory_i._003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._005_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i._108_  (.A(\efabless_subsystem.reduction_memory_i._005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].sena ));
 sky130_fd_sc_hd__or3_2 \efabless_subsystem.reduction_memory_i._109_  (.A(\efabless_subsystem.reduction_memory_i.g17.Z[4] ),
    .B(\efabless_subsystem.reduction_memory_i.g17.Z[6] ),
    .C(\efabless_subsystem.reduction_memory_i.g17.Z[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._006_ ));
 sky130_fd_sc_hd__or4b_2 \efabless_subsystem.reduction_memory_i._110_  (.A(\efabless_subsystem.reduction_memory_i.g17.Z[2] ),
    .B(\efabless_subsystem.reduction_memory_i.g17.Z[3] ),
    .C(\efabless_subsystem.reduction_memory_i.g17.Z[5] ),
    .D_N(\efabless_subsystem.reduction_memory_i.g17.Z[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._007_ ));
 sky130_fd_sc_hd__or4_2 \efabless_subsystem.reduction_memory_i._111_  (.A(\efabless_subsystem.reduction_memory_i.g17.Z[1] ),
    .B(\efabless_subsystem.reduction_memory_i.g17.Z[0] ),
    .C(\efabless_subsystem.reduction_memory_i._006_ ),
    .D(\efabless_subsystem.reduction_memory_i._007_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._008_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i._112_  (.A(\efabless_subsystem.reduction_memory_i._008_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.UNCONNECTED102 ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.reduction_memory_i._113_  (.A(\efabless_subsystem._223_ ),
    .B(\efabless_subsystem.UNCONNECTED102 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._009_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i._114_  (.A(\efabless_subsystem.reduction_memory_i._009_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_85_26.g1.data1 ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i._115_  (.A(\efabless_subsystem._223_ ),
    .B(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .C(\efabless_subsystem.UNCONNECTED102 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i._010_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i._116_  (.A(\efabless_subsystem.reduction_memory_i._010_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.reduction_memory_i._117_  (.A1(\efabless_subsystem.reduction_memory_i._000_ ),
    .A2(\efabless_subsystem.compute_controller_i.o_red_params_pop ),
    .B1(\efabless_subsystem.reduction_memory_i._003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._118_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._015_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._119_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._016_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._120_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._017_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._121_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._018_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._122_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._019_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._123_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._020_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._124_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._021_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._125_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._022_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._126_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._023_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._127_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._024_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._128_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._025_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._129_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._026_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._130_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._027_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._131_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._028_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._132_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._029_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._133_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._030_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._134_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._031_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._135_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._032_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._136_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._033_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._137_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._034_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._138_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._035_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._139_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._036_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._140_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._037_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._141_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.reduction_memory_i._038_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._142_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._039_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._143_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._040_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._144_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._041_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._145_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._042_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._146_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._043_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._147_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._044_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._148_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._045_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._149_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._046_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._150_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._047_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._151_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._048_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._152_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._049_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._153_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._050_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._154_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._051_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._155_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._052_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._156_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._053_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._157_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._054_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._158_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._055_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._159_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._056_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._160_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._057_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._161_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._058_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._162_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._059_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._163_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._060_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._164_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._061_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._165_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._062_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._166_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._063_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._167_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._064_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._168_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._065_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._169_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._066_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._170_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._067_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._171_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._068_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._172_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._069_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._173_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._070_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._174_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._071_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._175_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._072_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._176_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._073_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._177_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._074_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._178_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._075_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._179_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._076_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._180_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._077_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._181_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._078_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._182_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._079_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._183_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._080_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._184_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._081_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._185_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._082_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._186_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._083_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._187_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._084_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._188_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._085_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._189_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._086_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._190_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._087_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._191_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._088_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._192_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._089_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._193_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._090_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._194_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._091_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._195_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._092_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._196_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._093_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._197_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._094_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._198_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._095_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._199_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._096_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.reduction_memory_i._200_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.reduction_memory_i._097_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i.add_144_39._12_  (.A(\efabless_subsystem.reduction_memory_i._015_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .C(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.reduction_memory_i.add_144_39._13_  (.A1(\efabless_subsystem.reduction_memory_i._015_ ),
    .A2(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .B1(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_144_39._01_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i.add_144_39._14_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_144_39.Z[1] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.reduction_memory_i.add_144_39._15_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i.add_144_39._16_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_144_39._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i.add_144_39._17_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39._02_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_144_39.Z[2] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.reduction_memory_i.add_144_39._18_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._04_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.add_144_39._19_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_144_39._05_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.reduction_memory_i.add_144_39._20_  (.A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_144_39._02_ ),
    .B1(\efabless_subsystem.reduction_memory_i.add_144_39._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39.Z[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.reduction_memory_i.add_144_39._21_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_144_39.Z[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.reduction_memory_i.add_144_39._22_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .C(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .D(\efabless_subsystem.reduction_memory_i.add_144_39._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._06_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.reduction_memory_i.add_144_39._23_  (.A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .A3(\efabless_subsystem.reduction_memory_i.add_144_39._04_ ),
    .B1(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._07_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.reduction_memory_i.add_144_39._24_  (.A_N(\efabless_subsystem.reduction_memory_i.add_144_39._06_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.add_144_39._25_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39.Z[5] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i.add_144_39._26_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .C(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._09_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i.add_144_39._27_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._04_ ),
    .C(\efabless_subsystem.reduction_memory_i.add_144_39._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._10_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.reduction_memory_i.add_144_39._28_  (.A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_144_39._06_ ),
    .B1_N(\efabless_subsystem.reduction_memory_i.add_144_39._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39.Z[6] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.reduction_memory_i.add_144_39._29_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._00_ ),
    .C(\efabless_subsystem.reduction_memory_i.add_144_39._04_ ),
    .D(\efabless_subsystem.reduction_memory_i.add_144_39._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39._11_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.reduction_memory_i.add_144_39._30_  (.A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_144_39._10_ ),
    .B1_N(\efabless_subsystem.reduction_memory_i.add_144_39._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.add_144_39._31_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39.Z[8] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.add_144_39._32_  (.A(\efabless_subsystem.reduction_memory_i._015_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_144_39.Z[0] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i.add_149_37._12_  (.A(\efabless_subsystem.reduction_memory_i._016_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .C(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ));
 sky130_fd_sc_hd__a21oi_2 \efabless_subsystem.reduction_memory_i.add_149_37._13_  (.A1(\efabless_subsystem.reduction_memory_i._016_ ),
    .A2(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .B1(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_149_37._01_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i.add_149_37._14_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_149_37.Z[1] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.reduction_memory_i.add_149_37._15_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._02_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i.add_149_37._16_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_149_37._03_ ));
 sky130_fd_sc_hd__nor2_2 \efabless_subsystem.reduction_memory_i.add_149_37._17_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37._02_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._03_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_149_37.Z[2] ));
 sky130_fd_sc_hd__and2_2 \efabless_subsystem.reduction_memory_i.add_149_37._18_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._04_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.add_149_37._19_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_149_37._05_ ));
 sky130_fd_sc_hd__o21a_2 \efabless_subsystem.reduction_memory_i.add_149_37._20_  (.A1(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_149_37._02_ ),
    .B1(\efabless_subsystem.reduction_memory_i.add_149_37._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37.Z[3] ));
 sky130_fd_sc_hd__xnor2_2 \efabless_subsystem.reduction_memory_i.add_149_37._21_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.add_149_37.Z[4] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.reduction_memory_i.add_149_37._22_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .C(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .D(\efabless_subsystem.reduction_memory_i.add_149_37._04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._06_ ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.reduction_memory_i.add_149_37._23_  (.A1(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .A3(\efabless_subsystem.reduction_memory_i.add_149_37._04_ ),
    .B1(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._07_ ));
 sky130_fd_sc_hd__and2b_2 \efabless_subsystem.reduction_memory_i.add_149_37._24_  (.A_N(\efabless_subsystem.reduction_memory_i.add_149_37._06_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._07_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._08_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.add_149_37._25_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37._08_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37.Z[5] ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i.add_149_37._26_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .C(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._09_ ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.reduction_memory_i.add_149_37._27_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._04_ ),
    .C(\efabless_subsystem.reduction_memory_i.add_149_37._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._10_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.reduction_memory_i.add_149_37._28_  (.A1(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_149_37._06_ ),
    .B1_N(\efabless_subsystem.reduction_memory_i.add_149_37._10_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37.Z[6] ));
 sky130_fd_sc_hd__and4_2 \efabless_subsystem.reduction_memory_i.add_149_37._29_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._00_ ),
    .C(\efabless_subsystem.reduction_memory_i.add_149_37._04_ ),
    .D(\efabless_subsystem.reduction_memory_i.add_149_37._09_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37._11_ ));
 sky130_fd_sc_hd__o21ba_2 \efabless_subsystem.reduction_memory_i.add_149_37._30_  (.A1(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .A2(\efabless_subsystem.reduction_memory_i.add_149_37._10_ ),
    .B1_N(\efabless_subsystem.reduction_memory_i.add_149_37._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.add_149_37._31_  (.A(\efabless_subsystem.reduction_memory_i.add_149_37.A[8] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37._11_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37.Z[8] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.add_149_37._32_  (.A(\efabless_subsystem.reduction_memory_i._016_ ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.add_149_37.Z[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19._0_  (.A(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19._1_  (.A(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[0] ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._08_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._039_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._09_  (.A0(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.in_0 ),
    .A1(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].d ),
    .S(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].sena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._10_  (.A0(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._040_ ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._11_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.in_0 ),
    .Q_N(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0]._06_ ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._0_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[0] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._1_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[1] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._2_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[2] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._3_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._4_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[4] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._5_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._6_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[6] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._7_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g17._8_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g17.Z[8] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._0_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[0] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._1_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[1] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._2_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[2] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._3_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[3] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._4_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[4] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._5_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[5] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._6_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[6] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._7_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[7] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.reduction_memory_i.g18._8_  (.A(\efabless_subsystem.reduction_memory_i.add_144_39.A[8] ),
    .B(\efabless_subsystem.reduction_memory_i.add_149_37.A[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.g18.Z[8] ));
 sky130_sram_0kbytes_1rw1r_24x32_8 \efabless_subsystem.reduction_memory_i.mem241  (.csb0(\efabless_subsystem.reduction_memory_i.n_160 ),
    .csb1(\efabless_subsystem.reduction_memory_i.n_162 ),
    .web0(\efabless_subsystem.reduction_memory_i.n_161 ),
    .clk0(wb_clk_i),
    .clk1(wb_clk_i),
    .addr0({\efabless_subsystem.reduction_memory_i.memory_addr[4] ,
    \efabless_subsystem.reduction_memory_i.memory_addr[3] ,
    \efabless_subsystem.reduction_memory_i.memory_addr[2] ,
    \efabless_subsystem.reduction_memory_i.memory_addr[1] ,
    \efabless_subsystem.reduction_memory_i.memory_addr[0] }),
    .addr1({\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ,
    \efabless_subsystem.reduction_memory_i.add_149_37.A[3] ,
    \efabless_subsystem.reduction_memory_i.add_149_37.A[2] ,
    \efabless_subsystem.reduction_memory_i.add_149_37.A[1] ,
    \efabless_subsystem.reduction_memory_i.add_149_37.A[0] }),
    .din0({\efabless_subsystem.reduction_memory_i._042_ ,
    \efabless_subsystem.reduction_memory_i._041_ ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[21] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[20] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[19] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[18] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[17] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[16] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[15] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[14] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[13] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[12] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[11] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[10] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[9] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[8] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[7] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[6] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[5] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[4] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[3] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[2] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[1] ,
    \efabless_subsystem.reduction_memory_i.memory_wdata[0] }),
    .dout0({\efabless_subsystem.reduction_memory_i._014_ ,
    \efabless_subsystem.reduction_memory_i._013_ ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[21] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[20] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[19] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[18] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[17] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[16] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[15] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[14] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[13] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[12] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[11] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[10] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[9] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[8] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[7] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[6] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[5] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[4] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[3] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[2] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[1] ,
    \efabless_subsystem.mmap_interconnect_i.i_rmem_rdata[0] }),
    .dout1({\efabless_subsystem.reduction_memory_i._012_ ,
    \efabless_subsystem.reduction_memory_i._011_ ,
    \efabless_subsystem.compute_core_i.i_acc_sign ,
    \efabless_subsystem.compute_core_i.i_acc_shift[4] ,
    \efabless_subsystem.compute_core_i.i_acc_shift[3] ,
    \efabless_subsystem.compute_core_i.i_acc_shift[2] ,
    \efabless_subsystem.compute_core_i.i_acc_shift[1] ,
    \efabless_subsystem.compute_core_i.i_acc_shift[0] ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[15].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[14].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[13].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[12].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[11].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[10].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[9].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[8].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[7].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[6].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[5].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[4].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[3].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[2].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[1].d ,
    \efabless_subsystem.compute_controller_i.arr_red_cycles_q_reg[0].d }),
    .wmask0({\efabless_subsystem.reduction_memory_i.memory_wmask[2] ,
    \efabless_subsystem.reduction_memory_i.memory_wmask[1] ,
    \efabless_subsystem.reduction_memory_i.memory_wmask[0] }));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[21] ),
    .A1(\efabless_subsystem._222_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[21] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g10._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[12] ),
    .A1(\efabless_subsystem._213_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g10._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g10._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g10._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[12] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g11._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[11] ),
    .A1(\efabless_subsystem._212_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g11._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g11._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g11._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[11] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g12._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[10] ),
    .A1(\efabless_subsystem._211_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g12._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g12._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g12._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[10] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g13._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[9] ),
    .A1(\efabless_subsystem._210_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g13._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g13._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g13._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[9] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g14._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[8] ),
    .A1(\efabless_subsystem._209_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g14._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g14._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g14._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[8] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g15._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[7] ),
    .A1(\efabless_subsystem._208_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g15._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g15._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g15._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[7] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g16._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[6] ),
    .A1(\efabless_subsystem._207_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g16._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g16._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g16._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[6] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g17._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[5] ),
    .A1(\efabless_subsystem._206_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g17._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g17._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g17._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[5] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g18._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[4] ),
    .A1(\efabless_subsystem._205_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g18._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g18._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g18._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g19._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[3] ),
    .A1(\efabless_subsystem._204_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g19._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g19._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g19._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g2._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[20] ),
    .A1(\efabless_subsystem._221_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g2._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[20] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g20._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[2] ),
    .A1(\efabless_subsystem._203_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g20._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g20._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g20._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g21._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[1] ),
    .A1(\efabless_subsystem._202_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g21._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g21._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g21._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g22._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[0] ),
    .A1(\efabless_subsystem._201_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g22._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g22._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g22._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g3._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[19] ),
    .A1(\efabless_subsystem._220_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g3._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[19] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g4._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[18] ),
    .A1(\efabless_subsystem._219_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g4._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[18] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g5._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[17] ),
    .A1(\efabless_subsystem._218_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g5._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[17] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g6._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[16] ),
    .A1(\efabless_subsystem._217_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g6._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[16] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g7._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[15] ),
    .A1(\efabless_subsystem._216_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g7._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[15] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[14] ),
    .A1(\efabless_subsystem._215_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g8._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[14] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_82_26.g9._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wdata[13] ),
    .A1(\efabless_subsystem._214_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_82_26.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_82_26.g9._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_82_26.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wdata[13] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_83_26.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[16] ),
    .A1(\efabless_subsystem.reduction_memory_i._019_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_83_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_83_26.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_83_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wmask[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_83_26.g2._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[8] ),
    .A1(\efabless_subsystem.reduction_memory_i._018_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_83_26.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_83_26.g2._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_83_26.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wmask[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_83_26.g3._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_wmask[0] ),
    .A1(\efabless_subsystem.reduction_memory_i._017_ ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_83_26.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_83_26.g3._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_83_26.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wmask[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_84_26.g4._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[4] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_84_26.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_84_26.g4._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_84_26.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_addr[4] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_84_26.g5._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[3] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_84_26.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_84_26.g5._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_84_26.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_addr[3] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_84_26.g6._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[2] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_84_26.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_84_26.g6._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_84_26.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_addr[2] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_84_26.g7._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[1] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_84_26.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_84_26.g7._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_84_26.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_addr[1] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_84_26.g8._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.o_rmem_address[0] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_84_26.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_84_26.g8._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_84_26.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_addr[0] ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_85_26.g1._1_  (.A0(\efabless_subsystem.mmap_interconnect_i.mux_107_36.g1.z ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_85_26.g1.data1 ),
    .S(\efabless_subsystem.config_regs_i.mem_mode_q_reg.q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_85_26.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_85_26.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_85_26.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.memory_wren ));
 sky130_fd_sc_hd__a22o_2 \efabless_subsystem.reduction_memory_i.mux_fifo_state_103_19.g1._0_  (.A1(\efabless_subsystem.reduction_memory_i._020_ ),
    .A2(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[1] ),
    .B1(\efabless_subsystem.reduction_memory_i._043_ ),
    .B2(\efabless_subsystem.reduction_memory_i.ctl_fifo_state_103_19.out_0[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].d ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[8] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[7] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[6] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[5] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[4] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[3] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[2] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[1] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_rdptr_init[0] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g1._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[8] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[8] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g2._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[7] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g2._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g3._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[6] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g3._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g4._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[5] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g4._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g5._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[4] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g5._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g6._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[3] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g6._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g7._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[2] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g7._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g8._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[1] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g8._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g9._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_149_37.Z[0] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g9._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_148_22.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[8] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[7] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[6] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[5] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[4] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[3] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[2] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[1] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9._1_  (.A0(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9.data0 ),
    .A1(\efabless_subsystem.config_regs_i.o_rmem_fifo_wrptr_init[0] ),
    .S(\efabless_subsystem.config_regs_i.o_fifo_ptrs_set ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9.z ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g1._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[8] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[8] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g1._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g2._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[7] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g2._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g2._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g2._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g3._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[6] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g3._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g3._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g3._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g4._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[5] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g4._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g4._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g4._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g5._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[4] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g5._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g5._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g5._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g6._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[3] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g6._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g6._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g6._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g7._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[2] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g7._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g7._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g7._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g8._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[1] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g8._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g8._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g8._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8.data0 ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g9._1_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .A1(\efabless_subsystem.reduction_memory_i.add_144_39.Z[0] ),
    .S(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.ctl ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g9._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g9._2_  (.A(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_143_33.g9._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9.data0 ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._044_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g9.z ),
    .S(\efabless_subsystem.reduction_memory_i._021_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._045_ ),
    .S(\efabless_subsystem.reduction_memory_i._046_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[0] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._047_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g8.z ),
    .S(\efabless_subsystem.reduction_memory_i._022_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._048_ ),
    .S(\efabless_subsystem.reduction_memory_i._049_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[1] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._050_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g7.z ),
    .S(\efabless_subsystem.reduction_memory_i._023_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._051_ ),
    .S(\efabless_subsystem.reduction_memory_i._052_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[2] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._053_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g6.z ),
    .S(\efabless_subsystem.reduction_memory_i._024_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._054_ ),
    .S(\efabless_subsystem.reduction_memory_i._055_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[3] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._056_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g5.z ),
    .S(\efabless_subsystem.reduction_memory_i._025_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._057_ ),
    .S(\efabless_subsystem.reduction_memory_i._058_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[4] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._059_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g4.z ),
    .S(\efabless_subsystem.reduction_memory_i._026_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._060_ ),
    .S(\efabless_subsystem.reduction_memory_i._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[5] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g3.z ),
    .S(\efabless_subsystem.reduction_memory_i._027_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._063_ ),
    .S(\efabless_subsystem.reduction_memory_i._064_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[6] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._065_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g2.z ),
    .S(\efabless_subsystem.reduction_memory_i._028_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._066_ ),
    .S(\efabless_subsystem.reduction_memory_i._067_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[7] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._08_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._068_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_149_37.A[8] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_read_ptr_d_135_9.g1.z ),
    .S(\efabless_subsystem.reduction_memory_i._029_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._10_  (.A0(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._069_ ),
    .S(\efabless_subsystem.reduction_memory_i._070_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._11_  (.A(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_149_37.A[8] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.read_ptr_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._071_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g9.z ),
    .S(\efabless_subsystem.reduction_memory_i._030_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._072_ ),
    .S(\efabless_subsystem.reduction_memory_i._073_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[0] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[0]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._074_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g8.z ),
    .S(\efabless_subsystem.reduction_memory_i._031_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._075_ ),
    .S(\efabless_subsystem.reduction_memory_i._076_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[1] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[1]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._077_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g7.z ),
    .S(\efabless_subsystem.reduction_memory_i._032_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._078_ ),
    .S(\efabless_subsystem.reduction_memory_i._079_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[2] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[2]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._080_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g6.z ),
    .S(\efabless_subsystem.reduction_memory_i._033_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._081_ ),
    .S(\efabless_subsystem.reduction_memory_i._082_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[3] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[3]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._083_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g5.z ),
    .S(\efabless_subsystem.reduction_memory_i._034_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._084_ ),
    .S(\efabless_subsystem.reduction_memory_i._085_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[4] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[4]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._086_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g4.z ),
    .S(\efabless_subsystem.reduction_memory_i._035_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._087_ ),
    .S(\efabless_subsystem.reduction_memory_i._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[5] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[5]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._089_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g3.z ),
    .S(\efabless_subsystem.reduction_memory_i._036_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._090_ ),
    .S(\efabless_subsystem.reduction_memory_i._091_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[6] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[6]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._092_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g2.z ),
    .S(\efabless_subsystem.reduction_memory_i._037_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._093_ ),
    .S(\efabless_subsystem.reduction_memory_i._094_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[7] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[7]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._07_  (.A(\efabless_subsystem.reduction_memory_i.fifo_state_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._08_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._00_ ),
    .B(\efabless_subsystem.reduction_memory_i._095_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._09_  (.A0(\efabless_subsystem.reduction_memory_i.add_144_39.A[8] ),
    .A1(\efabless_subsystem.reduction_memory_i.mux_write_ptr_d_135_9.g1.z ),
    .S(\efabless_subsystem.reduction_memory_i._038_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._10_  (.A0(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._04_ ),
    .A1(\efabless_subsystem.reduction_memory_i._096_ ),
    .S(\efabless_subsystem.reduction_memory_i._097_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._11_  (.A(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._13_  (.CLK_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._02_ ),
    .D(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._03_ ),
    .RESET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._00_ ),
    .SET_B(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.reduction_memory_i.add_144_39.A[8] ),
    .Q_N(\efabless_subsystem.reduction_memory_i.write_ptr_q_reg[8]._06_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.wishbone_2mmap_i._008_  (.A(wb_rst_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0].aclr ));
 sky130_fd_sc_hd__and3_2 \efabless_subsystem.wishbone_2mmap_i._009_  (.A(wbs_stb_i),
    .B(wbs_cyc_i),
    .C(wbs_we_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i._000_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.wishbone_2mmap_i._010_  (.A(\efabless_subsystem.wishbone_2mmap_i._000_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wren ));
 sky130_fd_sc_hd__and3b_2 \efabless_subsystem.wishbone_2mmap_i._011_  (.A_N(wbs_we_i),
    .B(wbs_cyc_i),
    .C(wbs_stb_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i._001_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.wishbone_2mmap_i._012_  (.A(\efabless_subsystem.wishbone_2mmap_i._001_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_rden ));
 sky130_fd_sc_hd__a31o_2 \efabless_subsystem.wishbone_2mmap_i._013_  (.A1(wbs_stb_i),
    .A2(wbs_cyc_i),
    .A3(wbs_we_i),
    .B1(\efabless_subsystem.wishbone_2mmap_i.ack_delayed ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.wishbone_2mmap_i._014_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.wishbone_2mmap_i._002_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.wishbone_2mmap_i._015_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.wishbone_2mmap_i._003_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.wishbone_2mmap_i._016_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(\efabless_subsystem.wishbone_2mmap_i._004_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.wishbone_2mmap_i._017_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.wishbone_2mmap_i._005_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.wishbone_2mmap_i._018_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.wishbone_2mmap_i._006_ ));
 sky130_fd_sc_hd__conb_1 \efabless_subsystem.wishbone_2mmap_i._019_  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(\efabless_subsystem.wishbone_2mmap_i._007_ ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._022_  (.A(wbs_adr_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._023_  (.A(wbs_adr_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._024_  (.A(wbs_adr_i[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._025_  (.A(wbs_adr_i[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._026_  (.A(wbs_adr_i[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._027_  (.A(wbs_adr_i[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._028_  (.A(wbs_adr_i[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._029_  (.A(wbs_adr_i[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._030_  (.A(wbs_adr_i[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._031_  (.A(wbs_adr_i[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._032_  (.A(wbs_adr_i[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._033_  (.A(wbs_adr_i[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._034_  (.A(wbs_adr_i[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._035_  (.A(wbs_adr_i[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._036_  (.A(wbs_adr_i[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._037_  (.A(wbs_adr_i[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._038_  (.A(wbs_adr_i[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._039_  (.A(wbs_adr_i[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._040_  (.A(wbs_adr_i[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._041_  (.A(wbs_adr_i[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._042_  (.A(wbs_adr_i[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._043_  (.A(wbs_adr_i[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_address[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._052_  (.A(wbs_dat_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._053_  (.A(wbs_dat_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._054_  (.A(wbs_dat_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._055_  (.A(wbs_dat_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._056_  (.A(wbs_dat_i[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._057_  (.A(wbs_dat_i[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._058_  (.A(wbs_dat_i[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._059_  (.A(wbs_dat_i[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._060_  (.A(wbs_dat_i[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._061_  (.A(wbs_dat_i[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._062_  (.A(wbs_dat_i[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._063_  (.A(wbs_dat_i[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._064_  (.A(wbs_dat_i[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._065_  (.A(wbs_dat_i[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._066_  (.A(wbs_dat_i[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._067_  (.A(wbs_dat_i[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._068_  (.A(wbs_dat_i[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._069_  (.A(wbs_dat_i[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._070_  (.A(wbs_dat_i[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._071_  (.A(wbs_dat_i[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._072_  (.A(wbs_dat_i[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._073_  (.A(wbs_dat_i[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._074_  (.A(wbs_dat_i[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._075_  (.A(wbs_dat_i[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._076_  (.A(wbs_dat_i[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._077_  (.A(wbs_dat_i[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._078_  (.A(wbs_dat_i[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._079_  (.A(wbs_dat_i[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._080_  (.A(wbs_dat_i[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._081_  (.A(wbs_dat_i[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._082_  (.A(wbs_dat_i[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[30] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._083_  (.A(wbs_dat_i[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wdata[31] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._084_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[0] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._085_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[1] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._086_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[2] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._087_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[3] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._088_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[4] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._089_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[5] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._090_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[6] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._091_  (.A(wbs_sel_i[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[7] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._092_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[8] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._093_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[9] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._094_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[10] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._095_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[11] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._096_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[12] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._097_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[13] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._098_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[14] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._099_  (.A(wbs_sel_i[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[15] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._100_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[16] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._101_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[17] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._102_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[18] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._103_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[19] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._104_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[20] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._105_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[21] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._106_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[22] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._107_  (.A(wbs_sel_i[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[23] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._108_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[24] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._109_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[25] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._110_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[26] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._111_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[27] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._112_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[28] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._113_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[29] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._114_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[30] ));
 sky130_fd_sc_hd__buf_2 \efabless_subsystem.wishbone_2mmap_i._115_  (.A(wbs_sel_i[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.cpu_wmask[31] ));
 sky130_fd_sc_hd__xor2_2 \efabless_subsystem.wishbone_2mmap_i.add_88_47._0_  (.A(\efabless_subsystem.wishbone_2mmap_i._002_ ),
    .B(\efabless_subsystem.wishbone_2mmap_i.add_88_47.A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.add_88_47.Z ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._07_  (.A(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0].aclr ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._00_ ));
 sky130_fd_sc_hd__nand2_2 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._08_  (.A(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._00_ ),
    .B(\efabless_subsystem.wishbone_2mmap_i._005_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._01_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._09_  (.A0(\efabless_subsystem.wishbone_2mmap_i.add_88_47.A ),
    .A1(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0].d ),
    .S(\efabless_subsystem.wishbone_2mmap_i._003_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._04_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._10_  (.A0(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._04_ ),
    .A1(\efabless_subsystem.wishbone_2mmap_i._006_ ),
    .S(\efabless_subsystem.wishbone_2mmap_i.add_88_47.A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._05_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._11_  (.A(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._03_ ));
 sky130_fd_sc_hd__inv_2 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._12_  (.A(wb_clk_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._02_ ));
 sky130_fd_sc_hd__dfbbn_2 \efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._13_  (.CLK_N(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._02_ ),
    .D(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._03_ ),
    .RESET_B(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._00_ ),
    .SET_B(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._01_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\efabless_subsystem.wishbone_2mmap_i.add_88_47.A ),
    .Q_N(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0]._06_ ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.wishbone_2mmap_i.mux_ack_delayed_83_27.g1._1_  (.A0(\efabless_subsystem.wishbone_2mmap_i._007_ ),
    .A1(\efabless_subsystem.wishbone_2mmap_i._004_ ),
    .S(\efabless_subsystem.wishbone_2mmap_i.add_88_47.A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.mux_ack_delayed_83_27.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.wishbone_2mmap_i.mux_ack_delayed_83_27.g1._2_  (.A(\efabless_subsystem.wishbone_2mmap_i.mux_ack_delayed_83_27.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.ack_delayed ));
 sky130_fd_sc_hd__mux2_2 \efabless_subsystem.wishbone_2mmap_i.mux_latency_cnt_d_87_17.g1._1_  (.A0(\efabless_subsystem.wishbone_2mmap_i.add_88_47.A ),
    .A1(\efabless_subsystem.wishbone_2mmap_i.add_88_47.Z ),
    .S(\efabless_subsystem.cpu_rden ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.mux_latency_cnt_d_87_17.g1._0_ ));
 sky130_fd_sc_hd__buf_1 \efabless_subsystem.wishbone_2mmap_i.mux_latency_cnt_d_87_17.g1._2_  (.A(\efabless_subsystem.wishbone_2mmap_i.mux_latency_cnt_d_87_17.g1._0_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\efabless_subsystem.wishbone_2mmap_i.latency_cnt_q_reg[0].d ));
endmodule
